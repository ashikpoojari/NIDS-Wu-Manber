

module Wu_Manber_ShiftSelector
(
  input clk,
  input rst,
  input [1280-1:0] comp_shift_wire,
  output [5-1:0] shift_wire
);

  wire [5-1:0] shift_wire2561;
  assign shift_wire2561 = comp_shift_wire[4:0];
  wire [5-1:0] shift_wire2562;
  assign shift_wire2562 = comp_shift_wire[9:5];
  wire [5-1:0] shift_wire2563;
  assign shift_wire2563 = comp_shift_wire[14:10];
  wire [5-1:0] shift_wire2564;
  assign shift_wire2564 = comp_shift_wire[19:15];
  wire [5-1:0] shift_wire2565;
  assign shift_wire2565 = comp_shift_wire[24:20];
  wire [5-1:0] shift_wire2566;
  assign shift_wire2566 = comp_shift_wire[29:25];
  wire [5-1:0] shift_wire2567;
  assign shift_wire2567 = comp_shift_wire[34:30];
  wire [5-1:0] shift_wire2568;
  assign shift_wire2568 = comp_shift_wire[39:35];
  wire [5-1:0] shift_wire2569;
  assign shift_wire2569 = comp_shift_wire[44:40];
  wire [5-1:0] shift_wire2570;
  assign shift_wire2570 = comp_shift_wire[49:45];
  wire [5-1:0] shift_wire2571;
  assign shift_wire2571 = comp_shift_wire[54:50];
  wire [5-1:0] shift_wire2572;
  assign shift_wire2572 = comp_shift_wire[59:55];
  wire [5-1:0] shift_wire2573;
  assign shift_wire2573 = comp_shift_wire[64:60];
  wire [5-1:0] shift_wire2574;
  assign shift_wire2574 = comp_shift_wire[69:65];
  wire [5-1:0] shift_wire2575;
  assign shift_wire2575 = comp_shift_wire[74:70];
  wire [5-1:0] shift_wire2576;
  assign shift_wire2576 = comp_shift_wire[79:75];
  wire [5-1:0] shift_wire2577;
  assign shift_wire2577 = comp_shift_wire[84:80];
  wire [5-1:0] shift_wire2578;
  assign shift_wire2578 = comp_shift_wire[89:85];
  wire [5-1:0] shift_wire2579;
  assign shift_wire2579 = comp_shift_wire[94:90];
  wire [5-1:0] shift_wire2580;
  assign shift_wire2580 = comp_shift_wire[99:95];
  wire [5-1:0] shift_wire2581;
  assign shift_wire2581 = comp_shift_wire[104:100];
  wire [5-1:0] shift_wire2582;
  assign shift_wire2582 = comp_shift_wire[109:105];
  wire [5-1:0] shift_wire2583;
  assign shift_wire2583 = comp_shift_wire[114:110];
  wire [5-1:0] shift_wire2584;
  assign shift_wire2584 = comp_shift_wire[119:115];
  wire [5-1:0] shift_wire2585;
  assign shift_wire2585 = comp_shift_wire[124:120];
  wire [5-1:0] shift_wire2586;
  assign shift_wire2586 = comp_shift_wire[129:125];
  wire [5-1:0] shift_wire2587;
  assign shift_wire2587 = comp_shift_wire[134:130];
  wire [5-1:0] shift_wire2588;
  assign shift_wire2588 = comp_shift_wire[139:135];
  wire [5-1:0] shift_wire2589;
  assign shift_wire2589 = comp_shift_wire[144:140];
  wire [5-1:0] shift_wire2590;
  assign shift_wire2590 = comp_shift_wire[149:145];
  wire [5-1:0] shift_wire2591;
  assign shift_wire2591 = comp_shift_wire[154:150];
  wire [5-1:0] shift_wire2592;
  assign shift_wire2592 = comp_shift_wire[159:155];
  wire [5-1:0] shift_wire2593;
  assign shift_wire2593 = comp_shift_wire[164:160];
  wire [5-1:0] shift_wire2594;
  assign shift_wire2594 = comp_shift_wire[169:165];
  wire [5-1:0] shift_wire2595;
  assign shift_wire2595 = comp_shift_wire[174:170];
  wire [5-1:0] shift_wire2596;
  assign shift_wire2596 = comp_shift_wire[179:175];
  wire [5-1:0] shift_wire2597;
  assign shift_wire2597 = comp_shift_wire[184:180];
  wire [5-1:0] shift_wire2598;
  assign shift_wire2598 = comp_shift_wire[189:185];
  wire [5-1:0] shift_wire2599;
  assign shift_wire2599 = comp_shift_wire[194:190];
  wire [5-1:0] shift_wire2600;
  assign shift_wire2600 = comp_shift_wire[199:195];
  wire [5-1:0] shift_wire2601;
  assign shift_wire2601 = comp_shift_wire[204:200];
  wire [5-1:0] shift_wire2602;
  assign shift_wire2602 = comp_shift_wire[209:205];
  wire [5-1:0] shift_wire2603;
  assign shift_wire2603 = comp_shift_wire[214:210];
  wire [5-1:0] shift_wire2604;
  assign shift_wire2604 = comp_shift_wire[219:215];
  wire [5-1:0] shift_wire2605;
  assign shift_wire2605 = comp_shift_wire[224:220];
  wire [5-1:0] shift_wire2606;
  assign shift_wire2606 = comp_shift_wire[229:225];
  wire [5-1:0] shift_wire2607;
  assign shift_wire2607 = comp_shift_wire[234:230];
  wire [5-1:0] shift_wire2608;
  assign shift_wire2608 = comp_shift_wire[239:235];
  wire [5-1:0] shift_wire2609;
  assign shift_wire2609 = comp_shift_wire[244:240];
  wire [5-1:0] shift_wire2610;
  assign shift_wire2610 = comp_shift_wire[249:245];
  wire [5-1:0] shift_wire2611;
  assign shift_wire2611 = comp_shift_wire[254:250];
  wire [5-1:0] shift_wire2612;
  assign shift_wire2612 = comp_shift_wire[259:255];
  wire [5-1:0] shift_wire2613;
  assign shift_wire2613 = comp_shift_wire[264:260];
  wire [5-1:0] shift_wire2614;
  assign shift_wire2614 = comp_shift_wire[269:265];
  wire [5-1:0] shift_wire2615;
  assign shift_wire2615 = comp_shift_wire[274:270];
  wire [5-1:0] shift_wire2616;
  assign shift_wire2616 = comp_shift_wire[279:275];
  wire [5-1:0] shift_wire2617;
  assign shift_wire2617 = comp_shift_wire[284:280];
  wire [5-1:0] shift_wire2618;
  assign shift_wire2618 = comp_shift_wire[289:285];
  wire [5-1:0] shift_wire2619;
  assign shift_wire2619 = comp_shift_wire[294:290];
  wire [5-1:0] shift_wire2620;
  assign shift_wire2620 = comp_shift_wire[299:295];
  wire [5-1:0] shift_wire2621;
  assign shift_wire2621 = comp_shift_wire[304:300];
  wire [5-1:0] shift_wire2622;
  assign shift_wire2622 = comp_shift_wire[309:305];
  wire [5-1:0] shift_wire2623;
  assign shift_wire2623 = comp_shift_wire[314:310];
  wire [5-1:0] shift_wire2624;
  assign shift_wire2624 = comp_shift_wire[319:315];
  wire [5-1:0] shift_wire2625;
  assign shift_wire2625 = comp_shift_wire[324:320];
  wire [5-1:0] shift_wire2626;
  assign shift_wire2626 = comp_shift_wire[329:325];
  wire [5-1:0] shift_wire2627;
  assign shift_wire2627 = comp_shift_wire[334:330];
  wire [5-1:0] shift_wire2628;
  assign shift_wire2628 = comp_shift_wire[339:335];
  wire [5-1:0] shift_wire2629;
  assign shift_wire2629 = comp_shift_wire[344:340];
  wire [5-1:0] shift_wire2630;
  assign shift_wire2630 = comp_shift_wire[349:345];
  wire [5-1:0] shift_wire2631;
  assign shift_wire2631 = comp_shift_wire[354:350];
  wire [5-1:0] shift_wire2632;
  assign shift_wire2632 = comp_shift_wire[359:355];
  wire [5-1:0] shift_wire2633;
  assign shift_wire2633 = comp_shift_wire[364:360];
  wire [5-1:0] shift_wire2634;
  assign shift_wire2634 = comp_shift_wire[369:365];
  wire [5-1:0] shift_wire2635;
  assign shift_wire2635 = comp_shift_wire[374:370];
  wire [5-1:0] shift_wire2636;
  assign shift_wire2636 = comp_shift_wire[379:375];
  wire [5-1:0] shift_wire2637;
  assign shift_wire2637 = comp_shift_wire[384:380];
  wire [5-1:0] shift_wire2638;
  assign shift_wire2638 = comp_shift_wire[389:385];
  wire [5-1:0] shift_wire2639;
  assign shift_wire2639 = comp_shift_wire[394:390];
  wire [5-1:0] shift_wire2640;
  assign shift_wire2640 = comp_shift_wire[399:395];
  wire [5-1:0] shift_wire2641;
  assign shift_wire2641 = comp_shift_wire[404:400];
  wire [5-1:0] shift_wire2642;
  assign shift_wire2642 = comp_shift_wire[409:405];
  wire [5-1:0] shift_wire2643;
  assign shift_wire2643 = comp_shift_wire[414:410];
  wire [5-1:0] shift_wire2644;
  assign shift_wire2644 = comp_shift_wire[419:415];
  wire [5-1:0] shift_wire2645;
  assign shift_wire2645 = comp_shift_wire[424:420];
  wire [5-1:0] shift_wire2646;
  assign shift_wire2646 = comp_shift_wire[429:425];
  wire [5-1:0] shift_wire2647;
  assign shift_wire2647 = comp_shift_wire[434:430];
  wire [5-1:0] shift_wire2648;
  assign shift_wire2648 = comp_shift_wire[439:435];
  wire [5-1:0] shift_wire2649;
  assign shift_wire2649 = comp_shift_wire[444:440];
  wire [5-1:0] shift_wire2650;
  assign shift_wire2650 = comp_shift_wire[449:445];
  wire [5-1:0] shift_wire2651;
  assign shift_wire2651 = comp_shift_wire[454:450];
  wire [5-1:0] shift_wire2652;
  assign shift_wire2652 = comp_shift_wire[459:455];
  wire [5-1:0] shift_wire2653;
  assign shift_wire2653 = comp_shift_wire[464:460];
  wire [5-1:0] shift_wire2654;
  assign shift_wire2654 = comp_shift_wire[469:465];
  wire [5-1:0] shift_wire2655;
  assign shift_wire2655 = comp_shift_wire[474:470];
  wire [5-1:0] shift_wire2656;
  assign shift_wire2656 = comp_shift_wire[479:475];
  wire [5-1:0] shift_wire2657;
  assign shift_wire2657 = comp_shift_wire[484:480];
  wire [5-1:0] shift_wire2658;
  assign shift_wire2658 = comp_shift_wire[489:485];
  wire [5-1:0] shift_wire2659;
  assign shift_wire2659 = comp_shift_wire[494:490];
  wire [5-1:0] shift_wire2660;
  assign shift_wire2660 = comp_shift_wire[499:495];
  wire [5-1:0] shift_wire2661;
  assign shift_wire2661 = comp_shift_wire[504:500];
  wire [5-1:0] shift_wire2662;
  assign shift_wire2662 = comp_shift_wire[509:505];
  wire [5-1:0] shift_wire2663;
  assign shift_wire2663 = comp_shift_wire[514:510];
  wire [5-1:0] shift_wire2664;
  assign shift_wire2664 = comp_shift_wire[519:515];
  wire [5-1:0] shift_wire2665;
  assign shift_wire2665 = comp_shift_wire[524:520];
  wire [5-1:0] shift_wire2666;
  assign shift_wire2666 = comp_shift_wire[529:525];
  wire [5-1:0] shift_wire2667;
  assign shift_wire2667 = comp_shift_wire[534:530];
  wire [5-1:0] shift_wire2668;
  assign shift_wire2668 = comp_shift_wire[539:535];
  wire [5-1:0] shift_wire2669;
  assign shift_wire2669 = comp_shift_wire[544:540];
  wire [5-1:0] shift_wire2670;
  assign shift_wire2670 = comp_shift_wire[549:545];
  wire [5-1:0] shift_wire2671;
  assign shift_wire2671 = comp_shift_wire[554:550];
  wire [5-1:0] shift_wire2672;
  assign shift_wire2672 = comp_shift_wire[559:555];
  wire [5-1:0] shift_wire2673;
  assign shift_wire2673 = comp_shift_wire[564:560];
  wire [5-1:0] shift_wire2674;
  assign shift_wire2674 = comp_shift_wire[569:565];
  wire [5-1:0] shift_wire2675;
  assign shift_wire2675 = comp_shift_wire[574:570];
  wire [5-1:0] shift_wire2676;
  assign shift_wire2676 = comp_shift_wire[579:575];
  wire [5-1:0] shift_wire2677;
  assign shift_wire2677 = comp_shift_wire[584:580];
  wire [5-1:0] shift_wire2678;
  assign shift_wire2678 = comp_shift_wire[589:585];
  wire [5-1:0] shift_wire2679;
  assign shift_wire2679 = comp_shift_wire[594:590];
  wire [5-1:0] shift_wire2680;
  assign shift_wire2680 = comp_shift_wire[599:595];
  wire [5-1:0] shift_wire2681;
  assign shift_wire2681 = comp_shift_wire[604:600];
  wire [5-1:0] shift_wire2682;
  assign shift_wire2682 = comp_shift_wire[609:605];
  wire [5-1:0] shift_wire2683;
  assign shift_wire2683 = comp_shift_wire[614:610];
  wire [5-1:0] shift_wire2684;
  assign shift_wire2684 = comp_shift_wire[619:615];
  wire [5-1:0] shift_wire2685;
  assign shift_wire2685 = comp_shift_wire[624:620];
  wire [5-1:0] shift_wire2686;
  assign shift_wire2686 = comp_shift_wire[629:625];
  wire [5-1:0] shift_wire2687;
  assign shift_wire2687 = comp_shift_wire[634:630];
  wire [5-1:0] shift_wire2688;
  assign shift_wire2688 = comp_shift_wire[639:635];
  wire [5-1:0] shift_wire2689;
  assign shift_wire2689 = comp_shift_wire[644:640];
  wire [5-1:0] shift_wire2690;
  assign shift_wire2690 = comp_shift_wire[649:645];
  wire [5-1:0] shift_wire2691;
  assign shift_wire2691 = comp_shift_wire[654:650];
  wire [5-1:0] shift_wire2692;
  assign shift_wire2692 = comp_shift_wire[659:655];
  wire [5-1:0] shift_wire2693;
  assign shift_wire2693 = comp_shift_wire[664:660];
  wire [5-1:0] shift_wire2694;
  assign shift_wire2694 = comp_shift_wire[669:665];
  wire [5-1:0] shift_wire2695;
  assign shift_wire2695 = comp_shift_wire[674:670];
  wire [5-1:0] shift_wire2696;
  assign shift_wire2696 = comp_shift_wire[679:675];
  wire [5-1:0] shift_wire2697;
  assign shift_wire2697 = comp_shift_wire[684:680];
  wire [5-1:0] shift_wire2698;
  assign shift_wire2698 = comp_shift_wire[689:685];
  wire [5-1:0] shift_wire2699;
  assign shift_wire2699 = comp_shift_wire[694:690];
  wire [5-1:0] shift_wire2700;
  assign shift_wire2700 = comp_shift_wire[699:695];
  wire [5-1:0] shift_wire2701;
  assign shift_wire2701 = comp_shift_wire[704:700];
  wire [5-1:0] shift_wire2702;
  assign shift_wire2702 = comp_shift_wire[709:705];
  wire [5-1:0] shift_wire2703;
  assign shift_wire2703 = comp_shift_wire[714:710];
  wire [5-1:0] shift_wire2704;
  assign shift_wire2704 = comp_shift_wire[719:715];
  wire [5-1:0] shift_wire2705;
  assign shift_wire2705 = comp_shift_wire[724:720];
  wire [5-1:0] shift_wire2706;
  assign shift_wire2706 = comp_shift_wire[729:725];
  wire [5-1:0] shift_wire2707;
  assign shift_wire2707 = comp_shift_wire[734:730];
  wire [5-1:0] shift_wire2708;
  assign shift_wire2708 = comp_shift_wire[739:735];
  wire [5-1:0] shift_wire2709;
  assign shift_wire2709 = comp_shift_wire[744:740];
  wire [5-1:0] shift_wire2710;
  assign shift_wire2710 = comp_shift_wire[749:745];
  wire [5-1:0] shift_wire2711;
  assign shift_wire2711 = comp_shift_wire[754:750];
  wire [5-1:0] shift_wire2712;
  assign shift_wire2712 = comp_shift_wire[759:755];
  wire [5-1:0] shift_wire2713;
  assign shift_wire2713 = comp_shift_wire[764:760];
  wire [5-1:0] shift_wire2714;
  assign shift_wire2714 = comp_shift_wire[769:765];
  wire [5-1:0] shift_wire2715;
  assign shift_wire2715 = comp_shift_wire[774:770];
  wire [5-1:0] shift_wire2716;
  assign shift_wire2716 = comp_shift_wire[779:775];
  wire [5-1:0] shift_wire2717;
  assign shift_wire2717 = comp_shift_wire[784:780];
  wire [5-1:0] shift_wire2718;
  assign shift_wire2718 = comp_shift_wire[789:785];
  wire [5-1:0] shift_wire2719;
  assign shift_wire2719 = comp_shift_wire[794:790];
  wire [5-1:0] shift_wire2720;
  assign shift_wire2720 = comp_shift_wire[799:795];
  wire [5-1:0] shift_wire2721;
  assign shift_wire2721 = comp_shift_wire[804:800];
  wire [5-1:0] shift_wire2722;
  assign shift_wire2722 = comp_shift_wire[809:805];
  wire [5-1:0] shift_wire2723;
  assign shift_wire2723 = comp_shift_wire[814:810];
  wire [5-1:0] shift_wire2724;
  assign shift_wire2724 = comp_shift_wire[819:815];
  wire [5-1:0] shift_wire2725;
  assign shift_wire2725 = comp_shift_wire[824:820];
  wire [5-1:0] shift_wire2726;
  assign shift_wire2726 = comp_shift_wire[829:825];
  wire [5-1:0] shift_wire2727;
  assign shift_wire2727 = comp_shift_wire[834:830];
  wire [5-1:0] shift_wire2728;
  assign shift_wire2728 = comp_shift_wire[839:835];
  wire [5-1:0] shift_wire2729;
  assign shift_wire2729 = comp_shift_wire[844:840];
  wire [5-1:0] shift_wire2730;
  assign shift_wire2730 = comp_shift_wire[849:845];
  wire [5-1:0] shift_wire2731;
  assign shift_wire2731 = comp_shift_wire[854:850];
  wire [5-1:0] shift_wire2732;
  assign shift_wire2732 = comp_shift_wire[859:855];
  wire [5-1:0] shift_wire2733;
  assign shift_wire2733 = comp_shift_wire[864:860];
  wire [5-1:0] shift_wire2734;
  assign shift_wire2734 = comp_shift_wire[869:865];
  wire [5-1:0] shift_wire2735;
  assign shift_wire2735 = comp_shift_wire[874:870];
  wire [5-1:0] shift_wire2736;
  assign shift_wire2736 = comp_shift_wire[879:875];
  wire [5-1:0] shift_wire2737;
  assign shift_wire2737 = comp_shift_wire[884:880];
  wire [5-1:0] shift_wire2738;
  assign shift_wire2738 = comp_shift_wire[889:885];
  wire [5-1:0] shift_wire2739;
  assign shift_wire2739 = comp_shift_wire[894:890];
  wire [5-1:0] shift_wire2740;
  assign shift_wire2740 = comp_shift_wire[899:895];
  wire [5-1:0] shift_wire2741;
  assign shift_wire2741 = comp_shift_wire[904:900];
  wire [5-1:0] shift_wire2742;
  assign shift_wire2742 = comp_shift_wire[909:905];
  wire [5-1:0] shift_wire2743;
  assign shift_wire2743 = comp_shift_wire[914:910];
  wire [5-1:0] shift_wire2744;
  assign shift_wire2744 = comp_shift_wire[919:915];
  wire [5-1:0] shift_wire2745;
  assign shift_wire2745 = comp_shift_wire[924:920];
  wire [5-1:0] shift_wire2746;
  assign shift_wire2746 = comp_shift_wire[929:925];
  wire [5-1:0] shift_wire2747;
  assign shift_wire2747 = comp_shift_wire[934:930];
  wire [5-1:0] shift_wire2748;
  assign shift_wire2748 = comp_shift_wire[939:935];
  wire [5-1:0] shift_wire2749;
  assign shift_wire2749 = comp_shift_wire[944:940];
  wire [5-1:0] shift_wire2750;
  assign shift_wire2750 = comp_shift_wire[949:945];
  wire [5-1:0] shift_wire2751;
  assign shift_wire2751 = comp_shift_wire[954:950];
  wire [5-1:0] shift_wire2752;
  assign shift_wire2752 = comp_shift_wire[959:955];
  wire [5-1:0] shift_wire2753;
  assign shift_wire2753 = comp_shift_wire[964:960];
  wire [5-1:0] shift_wire2754;
  assign shift_wire2754 = comp_shift_wire[969:965];
  wire [5-1:0] shift_wire2755;
  assign shift_wire2755 = comp_shift_wire[974:970];
  wire [5-1:0] shift_wire2756;
  assign shift_wire2756 = comp_shift_wire[979:975];
  wire [5-1:0] shift_wire2757;
  assign shift_wire2757 = comp_shift_wire[984:980];
  wire [5-1:0] shift_wire2758;
  assign shift_wire2758 = comp_shift_wire[989:985];
  wire [5-1:0] shift_wire2759;
  assign shift_wire2759 = comp_shift_wire[994:990];
  wire [5-1:0] shift_wire2760;
  assign shift_wire2760 = comp_shift_wire[999:995];
  wire [5-1:0] shift_wire2761;
  assign shift_wire2761 = comp_shift_wire[1004:1000];
  wire [5-1:0] shift_wire2762;
  assign shift_wire2762 = comp_shift_wire[1009:1005];
  wire [5-1:0] shift_wire2763;
  assign shift_wire2763 = comp_shift_wire[1014:1010];
  wire [5-1:0] shift_wire2764;
  assign shift_wire2764 = comp_shift_wire[1019:1015];
  wire [5-1:0] shift_wire2765;
  assign shift_wire2765 = comp_shift_wire[1024:1020];
  wire [5-1:0] shift_wire2766;
  assign shift_wire2766 = comp_shift_wire[1029:1025];
  wire [5-1:0] shift_wire2767;
  assign shift_wire2767 = comp_shift_wire[1034:1030];
  wire [5-1:0] shift_wire2768;
  assign shift_wire2768 = comp_shift_wire[1039:1035];
  wire [5-1:0] shift_wire2769;
  assign shift_wire2769 = comp_shift_wire[1044:1040];
  wire [5-1:0] shift_wire2770;
  assign shift_wire2770 = comp_shift_wire[1049:1045];
  wire [5-1:0] shift_wire2771;
  assign shift_wire2771 = comp_shift_wire[1054:1050];
  wire [5-1:0] shift_wire2772;
  assign shift_wire2772 = comp_shift_wire[1059:1055];
  wire [5-1:0] shift_wire2773;
  assign shift_wire2773 = comp_shift_wire[1064:1060];
  wire [5-1:0] shift_wire2774;
  assign shift_wire2774 = comp_shift_wire[1069:1065];
  wire [5-1:0] shift_wire2775;
  assign shift_wire2775 = comp_shift_wire[1074:1070];
  wire [5-1:0] shift_wire2776;
  assign shift_wire2776 = comp_shift_wire[1079:1075];
  wire [5-1:0] shift_wire2777;
  assign shift_wire2777 = comp_shift_wire[1084:1080];
  wire [5-1:0] shift_wire2778;
  assign shift_wire2778 = comp_shift_wire[1089:1085];
  wire [5-1:0] shift_wire2779;
  assign shift_wire2779 = comp_shift_wire[1094:1090];
  wire [5-1:0] shift_wire2780;
  assign shift_wire2780 = comp_shift_wire[1099:1095];
  wire [5-1:0] shift_wire2781;
  assign shift_wire2781 = comp_shift_wire[1104:1100];
  wire [5-1:0] shift_wire2782;
  assign shift_wire2782 = comp_shift_wire[1109:1105];
  wire [5-1:0] shift_wire2783;
  assign shift_wire2783 = comp_shift_wire[1114:1110];
  wire [5-1:0] shift_wire2784;
  assign shift_wire2784 = comp_shift_wire[1119:1115];
  wire [5-1:0] shift_wire2785;
  assign shift_wire2785 = comp_shift_wire[1124:1120];
  wire [5-1:0] shift_wire2786;
  assign shift_wire2786 = comp_shift_wire[1129:1125];
  wire [5-1:0] shift_wire2787;
  assign shift_wire2787 = comp_shift_wire[1134:1130];
  wire [5-1:0] shift_wire2788;
  assign shift_wire2788 = comp_shift_wire[1139:1135];
  wire [5-1:0] shift_wire2789;
  assign shift_wire2789 = comp_shift_wire[1144:1140];
  wire [5-1:0] shift_wire2790;
  assign shift_wire2790 = comp_shift_wire[1149:1145];
  wire [5-1:0] shift_wire2791;
  assign shift_wire2791 = comp_shift_wire[1154:1150];
  wire [5-1:0] shift_wire2792;
  assign shift_wire2792 = comp_shift_wire[1159:1155];
  wire [5-1:0] shift_wire2793;
  assign shift_wire2793 = comp_shift_wire[1164:1160];
  wire [5-1:0] shift_wire2794;
  assign shift_wire2794 = comp_shift_wire[1169:1165];
  wire [5-1:0] shift_wire2795;
  assign shift_wire2795 = comp_shift_wire[1174:1170];
  wire [5-1:0] shift_wire2796;
  assign shift_wire2796 = comp_shift_wire[1179:1175];
  wire [5-1:0] shift_wire2797;
  assign shift_wire2797 = comp_shift_wire[1184:1180];
  wire [5-1:0] shift_wire2798;
  assign shift_wire2798 = comp_shift_wire[1189:1185];
  wire [5-1:0] shift_wire2799;
  assign shift_wire2799 = comp_shift_wire[1194:1190];
  wire [5-1:0] shift_wire2800;
  assign shift_wire2800 = comp_shift_wire[1199:1195];
  wire [5-1:0] shift_wire2801;
  assign shift_wire2801 = comp_shift_wire[1204:1200];
  wire [5-1:0] shift_wire2802;
  assign shift_wire2802 = comp_shift_wire[1209:1205];
  wire [5-1:0] shift_wire2803;
  assign shift_wire2803 = comp_shift_wire[1214:1210];
  wire [5-1:0] shift_wire2804;
  assign shift_wire2804 = comp_shift_wire[1219:1215];
  wire [5-1:0] shift_wire2805;
  assign shift_wire2805 = comp_shift_wire[1224:1220];
  wire [5-1:0] shift_wire2806;
  assign shift_wire2806 = comp_shift_wire[1229:1225];
  wire [5-1:0] shift_wire2807;
  assign shift_wire2807 = comp_shift_wire[1234:1230];
  wire [5-1:0] shift_wire2808;
  assign shift_wire2808 = comp_shift_wire[1239:1235];
  wire [5-1:0] shift_wire2809;
  assign shift_wire2809 = comp_shift_wire[1244:1240];
  wire [5-1:0] shift_wire2810;
  assign shift_wire2810 = comp_shift_wire[1249:1245];
  wire [5-1:0] shift_wire2811;
  assign shift_wire2811 = comp_shift_wire[1254:1250];
  wire [5-1:0] shift_wire2812;
  assign shift_wire2812 = comp_shift_wire[1259:1255];
  wire [5-1:0] shift_wire2813;
  assign shift_wire2813 = comp_shift_wire[1264:1260];
  wire [5-1:0] shift_wire2814;
  assign shift_wire2814 = comp_shift_wire[1269:1265];
  wire [5-1:0] shift_wire2815;
  assign shift_wire2815 = comp_shift_wire[1274:1270];
  wire [5-1:0] shift_wire2816;
  assign shift_wire2816 = comp_shift_wire[1279:1275];
  wire [5-1:0] shift_wire1281;

  muxaltb
  muxcmp1281
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2561),
    .b(shift_wire2562),
    .c(shift_wire1281)
  );

  wire [5-1:0] shift_wire1282;

  muxaltb
  muxcmp1282
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2563),
    .b(shift_wire2564),
    .c(shift_wire1282)
  );

  wire [5-1:0] shift_wire1283;

  muxaltb
  muxcmp1283
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2565),
    .b(shift_wire2566),
    .c(shift_wire1283)
  );

  wire [5-1:0] shift_wire1284;

  muxaltb
  muxcmp1284
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2567),
    .b(shift_wire2568),
    .c(shift_wire1284)
  );

  wire [5-1:0] shift_wire1285;

  muxaltb
  muxcmp1285
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2569),
    .b(shift_wire2570),
    .c(shift_wire1285)
  );

  wire [5-1:0] shift_wire1286;

  muxaltb
  muxcmp1286
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2571),
    .b(shift_wire2572),
    .c(shift_wire1286)
  );

  wire [5-1:0] shift_wire1287;

  muxaltb
  muxcmp1287
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2573),
    .b(shift_wire2574),
    .c(shift_wire1287)
  );

  wire [5-1:0] shift_wire1288;

  muxaltb
  muxcmp1288
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2575),
    .b(shift_wire2576),
    .c(shift_wire1288)
  );

  wire [5-1:0] shift_wire1289;

  muxaltb
  muxcmp1289
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2577),
    .b(shift_wire2578),
    .c(shift_wire1289)
  );

  wire [5-1:0] shift_wire1290;

  muxaltb
  muxcmp1290
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2579),
    .b(shift_wire2580),
    .c(shift_wire1290)
  );

  wire [5-1:0] shift_wire1291;

  muxaltb
  muxcmp1291
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2581),
    .b(shift_wire2582),
    .c(shift_wire1291)
  );

  wire [5-1:0] shift_wire1292;

  muxaltb
  muxcmp1292
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2583),
    .b(shift_wire2584),
    .c(shift_wire1292)
  );

  wire [5-1:0] shift_wire1293;

  muxaltb
  muxcmp1293
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2585),
    .b(shift_wire2586),
    .c(shift_wire1293)
  );

  wire [5-1:0] shift_wire1294;

  muxaltb
  muxcmp1294
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2587),
    .b(shift_wire2588),
    .c(shift_wire1294)
  );

  wire [5-1:0] shift_wire1295;

  muxaltb
  muxcmp1295
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2589),
    .b(shift_wire2590),
    .c(shift_wire1295)
  );

  wire [5-1:0] shift_wire1296;

  muxaltb
  muxcmp1296
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2591),
    .b(shift_wire2592),
    .c(shift_wire1296)
  );

  wire [5-1:0] shift_wire1297;

  muxaltb
  muxcmp1297
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2593),
    .b(shift_wire2594),
    .c(shift_wire1297)
  );

  wire [5-1:0] shift_wire1298;

  muxaltb
  muxcmp1298
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2595),
    .b(shift_wire2596),
    .c(shift_wire1298)
  );

  wire [5-1:0] shift_wire1299;

  muxaltb
  muxcmp1299
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2597),
    .b(shift_wire2598),
    .c(shift_wire1299)
  );

  wire [5-1:0] shift_wire1300;

  muxaltb
  muxcmp1300
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2599),
    .b(shift_wire2600),
    .c(shift_wire1300)
  );

  wire [5-1:0] shift_wire1301;

  muxaltb
  muxcmp1301
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2601),
    .b(shift_wire2602),
    .c(shift_wire1301)
  );

  wire [5-1:0] shift_wire1302;

  muxaltb
  muxcmp1302
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2603),
    .b(shift_wire2604),
    .c(shift_wire1302)
  );

  wire [5-1:0] shift_wire1303;

  muxaltb
  muxcmp1303
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2605),
    .b(shift_wire2606),
    .c(shift_wire1303)
  );

  wire [5-1:0] shift_wire1304;

  muxaltb
  muxcmp1304
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2607),
    .b(shift_wire2608),
    .c(shift_wire1304)
  );

  wire [5-1:0] shift_wire1305;

  muxaltb
  muxcmp1305
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2609),
    .b(shift_wire2610),
    .c(shift_wire1305)
  );

  wire [5-1:0] shift_wire1306;

  muxaltb
  muxcmp1306
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2611),
    .b(shift_wire2612),
    .c(shift_wire1306)
  );

  wire [5-1:0] shift_wire1307;

  muxaltb
  muxcmp1307
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2613),
    .b(shift_wire2614),
    .c(shift_wire1307)
  );

  wire [5-1:0] shift_wire1308;

  muxaltb
  muxcmp1308
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2615),
    .b(shift_wire2616),
    .c(shift_wire1308)
  );

  wire [5-1:0] shift_wire1309;

  muxaltb
  muxcmp1309
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2617),
    .b(shift_wire2618),
    .c(shift_wire1309)
  );

  wire [5-1:0] shift_wire1310;

  muxaltb
  muxcmp1310
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2619),
    .b(shift_wire2620),
    .c(shift_wire1310)
  );

  wire [5-1:0] shift_wire1311;

  muxaltb
  muxcmp1311
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2621),
    .b(shift_wire2622),
    .c(shift_wire1311)
  );

  wire [5-1:0] shift_wire1312;

  muxaltb
  muxcmp1312
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2623),
    .b(shift_wire2624),
    .c(shift_wire1312)
  );

  wire [5-1:0] shift_wire1313;

  muxaltb
  muxcmp1313
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2625),
    .b(shift_wire2626),
    .c(shift_wire1313)
  );

  wire [5-1:0] shift_wire1314;

  muxaltb
  muxcmp1314
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2627),
    .b(shift_wire2628),
    .c(shift_wire1314)
  );

  wire [5-1:0] shift_wire1315;

  muxaltb
  muxcmp1315
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2629),
    .b(shift_wire2630),
    .c(shift_wire1315)
  );

  wire [5-1:0] shift_wire1316;

  muxaltb
  muxcmp1316
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2631),
    .b(shift_wire2632),
    .c(shift_wire1316)
  );

  wire [5-1:0] shift_wire1317;

  muxaltb
  muxcmp1317
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2633),
    .b(shift_wire2634),
    .c(shift_wire1317)
  );

  wire [5-1:0] shift_wire1318;

  muxaltb
  muxcmp1318
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2635),
    .b(shift_wire2636),
    .c(shift_wire1318)
  );

  wire [5-1:0] shift_wire1319;

  muxaltb
  muxcmp1319
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2637),
    .b(shift_wire2638),
    .c(shift_wire1319)
  );

  wire [5-1:0] shift_wire1320;

  muxaltb
  muxcmp1320
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2639),
    .b(shift_wire2640),
    .c(shift_wire1320)
  );

  wire [5-1:0] shift_wire1321;

  muxaltb
  muxcmp1321
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2641),
    .b(shift_wire2642),
    .c(shift_wire1321)
  );

  wire [5-1:0] shift_wire1322;

  muxaltb
  muxcmp1322
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2643),
    .b(shift_wire2644),
    .c(shift_wire1322)
  );

  wire [5-1:0] shift_wire1323;

  muxaltb
  muxcmp1323
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2645),
    .b(shift_wire2646),
    .c(shift_wire1323)
  );

  wire [5-1:0] shift_wire1324;

  muxaltb
  muxcmp1324
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2647),
    .b(shift_wire2648),
    .c(shift_wire1324)
  );

  wire [5-1:0] shift_wire1325;

  muxaltb
  muxcmp1325
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2649),
    .b(shift_wire2650),
    .c(shift_wire1325)
  );

  wire [5-1:0] shift_wire1326;

  muxaltb
  muxcmp1326
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2651),
    .b(shift_wire2652),
    .c(shift_wire1326)
  );

  wire [5-1:0] shift_wire1327;

  muxaltb
  muxcmp1327
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2653),
    .b(shift_wire2654),
    .c(shift_wire1327)
  );

  wire [5-1:0] shift_wire1328;

  muxaltb
  muxcmp1328
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2655),
    .b(shift_wire2656),
    .c(shift_wire1328)
  );

  wire [5-1:0] shift_wire1329;

  muxaltb
  muxcmp1329
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2657),
    .b(shift_wire2658),
    .c(shift_wire1329)
  );

  wire [5-1:0] shift_wire1330;

  muxaltb
  muxcmp1330
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2659),
    .b(shift_wire2660),
    .c(shift_wire1330)
  );

  wire [5-1:0] shift_wire1331;

  muxaltb
  muxcmp1331
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2661),
    .b(shift_wire2662),
    .c(shift_wire1331)
  );

  wire [5-1:0] shift_wire1332;

  muxaltb
  muxcmp1332
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2663),
    .b(shift_wire2664),
    .c(shift_wire1332)
  );

  wire [5-1:0] shift_wire1333;

  muxaltb
  muxcmp1333
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2665),
    .b(shift_wire2666),
    .c(shift_wire1333)
  );

  wire [5-1:0] shift_wire1334;

  muxaltb
  muxcmp1334
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2667),
    .b(shift_wire2668),
    .c(shift_wire1334)
  );

  wire [5-1:0] shift_wire1335;

  muxaltb
  muxcmp1335
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2669),
    .b(shift_wire2670),
    .c(shift_wire1335)
  );

  wire [5-1:0] shift_wire1336;

  muxaltb
  muxcmp1336
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2671),
    .b(shift_wire2672),
    .c(shift_wire1336)
  );

  wire [5-1:0] shift_wire1337;

  muxaltb
  muxcmp1337
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2673),
    .b(shift_wire2674),
    .c(shift_wire1337)
  );

  wire [5-1:0] shift_wire1338;

  muxaltb
  muxcmp1338
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2675),
    .b(shift_wire2676),
    .c(shift_wire1338)
  );

  wire [5-1:0] shift_wire1339;

  muxaltb
  muxcmp1339
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2677),
    .b(shift_wire2678),
    .c(shift_wire1339)
  );

  wire [5-1:0] shift_wire1340;

  muxaltb
  muxcmp1340
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2679),
    .b(shift_wire2680),
    .c(shift_wire1340)
  );

  wire [5-1:0] shift_wire1341;

  muxaltb
  muxcmp1341
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2681),
    .b(shift_wire2682),
    .c(shift_wire1341)
  );

  wire [5-1:0] shift_wire1342;

  muxaltb
  muxcmp1342
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2683),
    .b(shift_wire2684),
    .c(shift_wire1342)
  );

  wire [5-1:0] shift_wire1343;

  muxaltb
  muxcmp1343
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2685),
    .b(shift_wire2686),
    .c(shift_wire1343)
  );

  wire [5-1:0] shift_wire1344;

  muxaltb
  muxcmp1344
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2687),
    .b(shift_wire2688),
    .c(shift_wire1344)
  );

  wire [5-1:0] shift_wire1345;

  muxaltb
  muxcmp1345
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2689),
    .b(shift_wire2690),
    .c(shift_wire1345)
  );

  wire [5-1:0] shift_wire1346;

  muxaltb
  muxcmp1346
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2691),
    .b(shift_wire2692),
    .c(shift_wire1346)
  );

  wire [5-1:0] shift_wire1347;

  muxaltb
  muxcmp1347
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2693),
    .b(shift_wire2694),
    .c(shift_wire1347)
  );

  wire [5-1:0] shift_wire1348;

  muxaltb
  muxcmp1348
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2695),
    .b(shift_wire2696),
    .c(shift_wire1348)
  );

  wire [5-1:0] shift_wire1349;

  muxaltb
  muxcmp1349
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2697),
    .b(shift_wire2698),
    .c(shift_wire1349)
  );

  wire [5-1:0] shift_wire1350;

  muxaltb
  muxcmp1350
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2699),
    .b(shift_wire2700),
    .c(shift_wire1350)
  );

  wire [5-1:0] shift_wire1351;

  muxaltb
  muxcmp1351
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2701),
    .b(shift_wire2702),
    .c(shift_wire1351)
  );

  wire [5-1:0] shift_wire1352;

  muxaltb
  muxcmp1352
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2703),
    .b(shift_wire2704),
    .c(shift_wire1352)
  );

  wire [5-1:0] shift_wire1353;

  muxaltb
  muxcmp1353
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2705),
    .b(shift_wire2706),
    .c(shift_wire1353)
  );

  wire [5-1:0] shift_wire1354;

  muxaltb
  muxcmp1354
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2707),
    .b(shift_wire2708),
    .c(shift_wire1354)
  );

  wire [5-1:0] shift_wire1355;

  muxaltb
  muxcmp1355
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2709),
    .b(shift_wire2710),
    .c(shift_wire1355)
  );

  wire [5-1:0] shift_wire1356;

  muxaltb
  muxcmp1356
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2711),
    .b(shift_wire2712),
    .c(shift_wire1356)
  );

  wire [5-1:0] shift_wire1357;

  muxaltb
  muxcmp1357
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2713),
    .b(shift_wire2714),
    .c(shift_wire1357)
  );

  wire [5-1:0] shift_wire1358;

  muxaltb
  muxcmp1358
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2715),
    .b(shift_wire2716),
    .c(shift_wire1358)
  );

  wire [5-1:0] shift_wire1359;

  muxaltb
  muxcmp1359
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2717),
    .b(shift_wire2718),
    .c(shift_wire1359)
  );

  wire [5-1:0] shift_wire1360;

  muxaltb
  muxcmp1360
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2719),
    .b(shift_wire2720),
    .c(shift_wire1360)
  );

  wire [5-1:0] shift_wire1361;

  muxaltb
  muxcmp1361
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2721),
    .b(shift_wire2722),
    .c(shift_wire1361)
  );

  wire [5-1:0] shift_wire1362;

  muxaltb
  muxcmp1362
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2723),
    .b(shift_wire2724),
    .c(shift_wire1362)
  );

  wire [5-1:0] shift_wire1363;

  muxaltb
  muxcmp1363
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2725),
    .b(shift_wire2726),
    .c(shift_wire1363)
  );

  wire [5-1:0] shift_wire1364;

  muxaltb
  muxcmp1364
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2727),
    .b(shift_wire2728),
    .c(shift_wire1364)
  );

  wire [5-1:0] shift_wire1365;

  muxaltb
  muxcmp1365
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2729),
    .b(shift_wire2730),
    .c(shift_wire1365)
  );

  wire [5-1:0] shift_wire1366;

  muxaltb
  muxcmp1366
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2731),
    .b(shift_wire2732),
    .c(shift_wire1366)
  );

  wire [5-1:0] shift_wire1367;

  muxaltb
  muxcmp1367
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2733),
    .b(shift_wire2734),
    .c(shift_wire1367)
  );

  wire [5-1:0] shift_wire1368;

  muxaltb
  muxcmp1368
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2735),
    .b(shift_wire2736),
    .c(shift_wire1368)
  );

  wire [5-1:0] shift_wire1369;

  muxaltb
  muxcmp1369
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2737),
    .b(shift_wire2738),
    .c(shift_wire1369)
  );

  wire [5-1:0] shift_wire1370;

  muxaltb
  muxcmp1370
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2739),
    .b(shift_wire2740),
    .c(shift_wire1370)
  );

  wire [5-1:0] shift_wire1371;

  muxaltb
  muxcmp1371
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2741),
    .b(shift_wire2742),
    .c(shift_wire1371)
  );

  wire [5-1:0] shift_wire1372;

  muxaltb
  muxcmp1372
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2743),
    .b(shift_wire2744),
    .c(shift_wire1372)
  );

  wire [5-1:0] shift_wire1373;

  muxaltb
  muxcmp1373
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2745),
    .b(shift_wire2746),
    .c(shift_wire1373)
  );

  wire [5-1:0] shift_wire1374;

  muxaltb
  muxcmp1374
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2747),
    .b(shift_wire2748),
    .c(shift_wire1374)
  );

  wire [5-1:0] shift_wire1375;

  muxaltb
  muxcmp1375
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2749),
    .b(shift_wire2750),
    .c(shift_wire1375)
  );

  wire [5-1:0] shift_wire1376;

  muxaltb
  muxcmp1376
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2751),
    .b(shift_wire2752),
    .c(shift_wire1376)
  );

  wire [5-1:0] shift_wire1377;

  muxaltb
  muxcmp1377
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2753),
    .b(shift_wire2754),
    .c(shift_wire1377)
  );

  wire [5-1:0] shift_wire1378;

  muxaltb
  muxcmp1378
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2755),
    .b(shift_wire2756),
    .c(shift_wire1378)
  );

  wire [5-1:0] shift_wire1379;

  muxaltb
  muxcmp1379
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2757),
    .b(shift_wire2758),
    .c(shift_wire1379)
  );

  wire [5-1:0] shift_wire1380;

  muxaltb
  muxcmp1380
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2759),
    .b(shift_wire2760),
    .c(shift_wire1380)
  );

  wire [5-1:0] shift_wire1381;

  muxaltb
  muxcmp1381
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2761),
    .b(shift_wire2762),
    .c(shift_wire1381)
  );

  wire [5-1:0] shift_wire1382;

  muxaltb
  muxcmp1382
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2763),
    .b(shift_wire2764),
    .c(shift_wire1382)
  );

  wire [5-1:0] shift_wire1383;

  muxaltb
  muxcmp1383
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2765),
    .b(shift_wire2766),
    .c(shift_wire1383)
  );

  wire [5-1:0] shift_wire1384;

  muxaltb
  muxcmp1384
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2767),
    .b(shift_wire2768),
    .c(shift_wire1384)
  );

  wire [5-1:0] shift_wire1385;

  muxaltb
  muxcmp1385
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2769),
    .b(shift_wire2770),
    .c(shift_wire1385)
  );

  wire [5-1:0] shift_wire1386;

  muxaltb
  muxcmp1386
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2771),
    .b(shift_wire2772),
    .c(shift_wire1386)
  );

  wire [5-1:0] shift_wire1387;

  muxaltb
  muxcmp1387
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2773),
    .b(shift_wire2774),
    .c(shift_wire1387)
  );

  wire [5-1:0] shift_wire1388;

  muxaltb
  muxcmp1388
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2775),
    .b(shift_wire2776),
    .c(shift_wire1388)
  );

  wire [5-1:0] shift_wire1389;

  muxaltb
  muxcmp1389
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2777),
    .b(shift_wire2778),
    .c(shift_wire1389)
  );

  wire [5-1:0] shift_wire1390;

  muxaltb
  muxcmp1390
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2779),
    .b(shift_wire2780),
    .c(shift_wire1390)
  );

  wire [5-1:0] shift_wire1391;

  muxaltb
  muxcmp1391
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2781),
    .b(shift_wire2782),
    .c(shift_wire1391)
  );

  wire [5-1:0] shift_wire1392;

  muxaltb
  muxcmp1392
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2783),
    .b(shift_wire2784),
    .c(shift_wire1392)
  );

  wire [5-1:0] shift_wire1393;

  muxaltb
  muxcmp1393
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2785),
    .b(shift_wire2786),
    .c(shift_wire1393)
  );

  wire [5-1:0] shift_wire1394;

  muxaltb
  muxcmp1394
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2787),
    .b(shift_wire2788),
    .c(shift_wire1394)
  );

  wire [5-1:0] shift_wire1395;

  muxaltb
  muxcmp1395
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2789),
    .b(shift_wire2790),
    .c(shift_wire1395)
  );

  wire [5-1:0] shift_wire1396;

  muxaltb
  muxcmp1396
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2791),
    .b(shift_wire2792),
    .c(shift_wire1396)
  );

  wire [5-1:0] shift_wire1397;

  muxaltb
  muxcmp1397
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2793),
    .b(shift_wire2794),
    .c(shift_wire1397)
  );

  wire [5-1:0] shift_wire1398;

  muxaltb
  muxcmp1398
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2795),
    .b(shift_wire2796),
    .c(shift_wire1398)
  );

  wire [5-1:0] shift_wire1399;

  muxaltb
  muxcmp1399
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2797),
    .b(shift_wire2798),
    .c(shift_wire1399)
  );

  wire [5-1:0] shift_wire1400;

  muxaltb
  muxcmp1400
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2799),
    .b(shift_wire2800),
    .c(shift_wire1400)
  );

  wire [5-1:0] shift_wire1401;

  muxaltb
  muxcmp1401
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2801),
    .b(shift_wire2802),
    .c(shift_wire1401)
  );

  wire [5-1:0] shift_wire1402;

  muxaltb
  muxcmp1402
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2803),
    .b(shift_wire2804),
    .c(shift_wire1402)
  );

  wire [5-1:0] shift_wire1403;

  muxaltb
  muxcmp1403
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2805),
    .b(shift_wire2806),
    .c(shift_wire1403)
  );

  wire [5-1:0] shift_wire1404;

  muxaltb
  muxcmp1404
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2807),
    .b(shift_wire2808),
    .c(shift_wire1404)
  );

  wire [5-1:0] shift_wire1405;

  muxaltb
  muxcmp1405
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2809),
    .b(shift_wire2810),
    .c(shift_wire1405)
  );

  wire [5-1:0] shift_wire1406;

  muxaltb
  muxcmp1406
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2811),
    .b(shift_wire2812),
    .c(shift_wire1406)
  );

  wire [5-1:0] shift_wire1407;

  muxaltb
  muxcmp1407
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2813),
    .b(shift_wire2814),
    .c(shift_wire1407)
  );

  wire [5-1:0] shift_wire1408;

  muxaltb
  muxcmp1408
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire2815),
    .b(shift_wire2816),
    .c(shift_wire1408)
  );

  wire [5-1:0] shift_wire641;

  muxaltb
  muxcmp641
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1281),
    .b(shift_wire1282),
    .c(shift_wire641)
  );

  wire [5-1:0] shift_wire642;

  muxaltb
  muxcmp642
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1283),
    .b(shift_wire1284),
    .c(shift_wire642)
  );

  wire [5-1:0] shift_wire643;

  muxaltb
  muxcmp643
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1285),
    .b(shift_wire1286),
    .c(shift_wire643)
  );

  wire [5-1:0] shift_wire644;

  muxaltb
  muxcmp644
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1287),
    .b(shift_wire1288),
    .c(shift_wire644)
  );

  wire [5-1:0] shift_wire645;

  muxaltb
  muxcmp645
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1289),
    .b(shift_wire1290),
    .c(shift_wire645)
  );

  wire [5-1:0] shift_wire646;

  muxaltb
  muxcmp646
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1291),
    .b(shift_wire1292),
    .c(shift_wire646)
  );

  wire [5-1:0] shift_wire647;

  muxaltb
  muxcmp647
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1293),
    .b(shift_wire1294),
    .c(shift_wire647)
  );

  wire [5-1:0] shift_wire648;

  muxaltb
  muxcmp648
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1295),
    .b(shift_wire1296),
    .c(shift_wire648)
  );

  wire [5-1:0] shift_wire649;

  muxaltb
  muxcmp649
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1297),
    .b(shift_wire1298),
    .c(shift_wire649)
  );

  wire [5-1:0] shift_wire650;

  muxaltb
  muxcmp650
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1299),
    .b(shift_wire1300),
    .c(shift_wire650)
  );

  wire [5-1:0] shift_wire651;

  muxaltb
  muxcmp651
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1301),
    .b(shift_wire1302),
    .c(shift_wire651)
  );

  wire [5-1:0] shift_wire652;

  muxaltb
  muxcmp652
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1303),
    .b(shift_wire1304),
    .c(shift_wire652)
  );

  wire [5-1:0] shift_wire653;

  muxaltb
  muxcmp653
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1305),
    .b(shift_wire1306),
    .c(shift_wire653)
  );

  wire [5-1:0] shift_wire654;

  muxaltb
  muxcmp654
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1307),
    .b(shift_wire1308),
    .c(shift_wire654)
  );

  wire [5-1:0] shift_wire655;

  muxaltb
  muxcmp655
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1309),
    .b(shift_wire1310),
    .c(shift_wire655)
  );

  wire [5-1:0] shift_wire656;

  muxaltb
  muxcmp656
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1311),
    .b(shift_wire1312),
    .c(shift_wire656)
  );

  wire [5-1:0] shift_wire657;

  muxaltb
  muxcmp657
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1313),
    .b(shift_wire1314),
    .c(shift_wire657)
  );

  wire [5-1:0] shift_wire658;

  muxaltb
  muxcmp658
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1315),
    .b(shift_wire1316),
    .c(shift_wire658)
  );

  wire [5-1:0] shift_wire659;

  muxaltb
  muxcmp659
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1317),
    .b(shift_wire1318),
    .c(shift_wire659)
  );

  wire [5-1:0] shift_wire660;

  muxaltb
  muxcmp660
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1319),
    .b(shift_wire1320),
    .c(shift_wire660)
  );

  wire [5-1:0] shift_wire661;

  muxaltb
  muxcmp661
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1321),
    .b(shift_wire1322),
    .c(shift_wire661)
  );

  wire [5-1:0] shift_wire662;

  muxaltb
  muxcmp662
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1323),
    .b(shift_wire1324),
    .c(shift_wire662)
  );

  wire [5-1:0] shift_wire663;

  muxaltb
  muxcmp663
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1325),
    .b(shift_wire1326),
    .c(shift_wire663)
  );

  wire [5-1:0] shift_wire664;

  muxaltb
  muxcmp664
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1327),
    .b(shift_wire1328),
    .c(shift_wire664)
  );

  wire [5-1:0] shift_wire665;

  muxaltb
  muxcmp665
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1329),
    .b(shift_wire1330),
    .c(shift_wire665)
  );

  wire [5-1:0] shift_wire666;

  muxaltb
  muxcmp666
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1331),
    .b(shift_wire1332),
    .c(shift_wire666)
  );

  wire [5-1:0] shift_wire667;

  muxaltb
  muxcmp667
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1333),
    .b(shift_wire1334),
    .c(shift_wire667)
  );

  wire [5-1:0] shift_wire668;

  muxaltb
  muxcmp668
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1335),
    .b(shift_wire1336),
    .c(shift_wire668)
  );

  wire [5-1:0] shift_wire669;

  muxaltb
  muxcmp669
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1337),
    .b(shift_wire1338),
    .c(shift_wire669)
  );

  wire [5-1:0] shift_wire670;

  muxaltb
  muxcmp670
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1339),
    .b(shift_wire1340),
    .c(shift_wire670)
  );

  wire [5-1:0] shift_wire671;

  muxaltb
  muxcmp671
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1341),
    .b(shift_wire1342),
    .c(shift_wire671)
  );

  wire [5-1:0] shift_wire672;

  muxaltb
  muxcmp672
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1343),
    .b(shift_wire1344),
    .c(shift_wire672)
  );

  wire [5-1:0] shift_wire673;

  muxaltb
  muxcmp673
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1345),
    .b(shift_wire1346),
    .c(shift_wire673)
  );

  wire [5-1:0] shift_wire674;

  muxaltb
  muxcmp674
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1347),
    .b(shift_wire1348),
    .c(shift_wire674)
  );

  wire [5-1:0] shift_wire675;

  muxaltb
  muxcmp675
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1349),
    .b(shift_wire1350),
    .c(shift_wire675)
  );

  wire [5-1:0] shift_wire676;

  muxaltb
  muxcmp676
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1351),
    .b(shift_wire1352),
    .c(shift_wire676)
  );

  wire [5-1:0] shift_wire677;

  muxaltb
  muxcmp677
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1353),
    .b(shift_wire1354),
    .c(shift_wire677)
  );

  wire [5-1:0] shift_wire678;

  muxaltb
  muxcmp678
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1355),
    .b(shift_wire1356),
    .c(shift_wire678)
  );

  wire [5-1:0] shift_wire679;

  muxaltb
  muxcmp679
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1357),
    .b(shift_wire1358),
    .c(shift_wire679)
  );

  wire [5-1:0] shift_wire680;

  muxaltb
  muxcmp680
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1359),
    .b(shift_wire1360),
    .c(shift_wire680)
  );

  wire [5-1:0] shift_wire681;

  muxaltb
  muxcmp681
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1361),
    .b(shift_wire1362),
    .c(shift_wire681)
  );

  wire [5-1:0] shift_wire682;

  muxaltb
  muxcmp682
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1363),
    .b(shift_wire1364),
    .c(shift_wire682)
  );

  wire [5-1:0] shift_wire683;

  muxaltb
  muxcmp683
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1365),
    .b(shift_wire1366),
    .c(shift_wire683)
  );

  wire [5-1:0] shift_wire684;

  muxaltb
  muxcmp684
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1367),
    .b(shift_wire1368),
    .c(shift_wire684)
  );

  wire [5-1:0] shift_wire685;

  muxaltb
  muxcmp685
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1369),
    .b(shift_wire1370),
    .c(shift_wire685)
  );

  wire [5-1:0] shift_wire686;

  muxaltb
  muxcmp686
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1371),
    .b(shift_wire1372),
    .c(shift_wire686)
  );

  wire [5-1:0] shift_wire687;

  muxaltb
  muxcmp687
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1373),
    .b(shift_wire1374),
    .c(shift_wire687)
  );

  wire [5-1:0] shift_wire688;

  muxaltb
  muxcmp688
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1375),
    .b(shift_wire1376),
    .c(shift_wire688)
  );

  wire [5-1:0] shift_wire689;

  muxaltb
  muxcmp689
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1377),
    .b(shift_wire1378),
    .c(shift_wire689)
  );

  wire [5-1:0] shift_wire690;

  muxaltb
  muxcmp690
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1379),
    .b(shift_wire1380),
    .c(shift_wire690)
  );

  wire [5-1:0] shift_wire691;

  muxaltb
  muxcmp691
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1381),
    .b(shift_wire1382),
    .c(shift_wire691)
  );

  wire [5-1:0] shift_wire692;

  muxaltb
  muxcmp692
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1383),
    .b(shift_wire1384),
    .c(shift_wire692)
  );

  wire [5-1:0] shift_wire693;

  muxaltb
  muxcmp693
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1385),
    .b(shift_wire1386),
    .c(shift_wire693)
  );

  wire [5-1:0] shift_wire694;

  muxaltb
  muxcmp694
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1387),
    .b(shift_wire1388),
    .c(shift_wire694)
  );

  wire [5-1:0] shift_wire695;

  muxaltb
  muxcmp695
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1389),
    .b(shift_wire1390),
    .c(shift_wire695)
  );

  wire [5-1:0] shift_wire696;

  muxaltb
  muxcmp696
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1391),
    .b(shift_wire1392),
    .c(shift_wire696)
  );

  wire [5-1:0] shift_wire697;

  muxaltb
  muxcmp697
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1393),
    .b(shift_wire1394),
    .c(shift_wire697)
  );

  wire [5-1:0] shift_wire698;

  muxaltb
  muxcmp698
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1395),
    .b(shift_wire1396),
    .c(shift_wire698)
  );

  wire [5-1:0] shift_wire699;

  muxaltb
  muxcmp699
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1397),
    .b(shift_wire1398),
    .c(shift_wire699)
  );

  wire [5-1:0] shift_wire700;

  muxaltb
  muxcmp700
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1399),
    .b(shift_wire1400),
    .c(shift_wire700)
  );

  wire [5-1:0] shift_wire701;

  muxaltb
  muxcmp701
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1401),
    .b(shift_wire1402),
    .c(shift_wire701)
  );

  wire [5-1:0] shift_wire702;

  muxaltb
  muxcmp702
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1403),
    .b(shift_wire1404),
    .c(shift_wire702)
  );

  wire [5-1:0] shift_wire703;

  muxaltb
  muxcmp703
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1405),
    .b(shift_wire1406),
    .c(shift_wire703)
  );

  wire [5-1:0] shift_wire704;

  muxaltb
  muxcmp704
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire1407),
    .b(shift_wire1408),
    .c(shift_wire704)
  );

  wire [5-1:0] shift_wire321;

  muxaltb
  muxcmp321
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire641),
    .b(shift_wire642),
    .c(shift_wire321)
  );

  wire [5-1:0] shift_wire322;

  muxaltb
  muxcmp322
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire643),
    .b(shift_wire644),
    .c(shift_wire322)
  );

  wire [5-1:0] shift_wire323;

  muxaltb
  muxcmp323
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire645),
    .b(shift_wire646),
    .c(shift_wire323)
  );

  wire [5-1:0] shift_wire324;

  muxaltb
  muxcmp324
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire647),
    .b(shift_wire648),
    .c(shift_wire324)
  );

  wire [5-1:0] shift_wire325;

  muxaltb
  muxcmp325
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire649),
    .b(shift_wire650),
    .c(shift_wire325)
  );

  wire [5-1:0] shift_wire326;

  muxaltb
  muxcmp326
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire651),
    .b(shift_wire652),
    .c(shift_wire326)
  );

  wire [5-1:0] shift_wire327;

  muxaltb
  muxcmp327
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire653),
    .b(shift_wire654),
    .c(shift_wire327)
  );

  wire [5-1:0] shift_wire328;

  muxaltb
  muxcmp328
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire655),
    .b(shift_wire656),
    .c(shift_wire328)
  );

  wire [5-1:0] shift_wire329;

  muxaltb
  muxcmp329
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire657),
    .b(shift_wire658),
    .c(shift_wire329)
  );

  wire [5-1:0] shift_wire330;

  muxaltb
  muxcmp330
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire659),
    .b(shift_wire660),
    .c(shift_wire330)
  );

  wire [5-1:0] shift_wire331;

  muxaltb
  muxcmp331
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire661),
    .b(shift_wire662),
    .c(shift_wire331)
  );

  wire [5-1:0] shift_wire332;

  muxaltb
  muxcmp332
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire663),
    .b(shift_wire664),
    .c(shift_wire332)
  );

  wire [5-1:0] shift_wire333;

  muxaltb
  muxcmp333
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire665),
    .b(shift_wire666),
    .c(shift_wire333)
  );

  wire [5-1:0] shift_wire334;

  muxaltb
  muxcmp334
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire667),
    .b(shift_wire668),
    .c(shift_wire334)
  );

  wire [5-1:0] shift_wire335;

  muxaltb
  muxcmp335
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire669),
    .b(shift_wire670),
    .c(shift_wire335)
  );

  wire [5-1:0] shift_wire336;

  muxaltb
  muxcmp336
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire671),
    .b(shift_wire672),
    .c(shift_wire336)
  );

  wire [5-1:0] shift_wire337;

  muxaltb
  muxcmp337
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire673),
    .b(shift_wire674),
    .c(shift_wire337)
  );

  wire [5-1:0] shift_wire338;

  muxaltb
  muxcmp338
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire675),
    .b(shift_wire676),
    .c(shift_wire338)
  );

  wire [5-1:0] shift_wire339;

  muxaltb
  muxcmp339
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire677),
    .b(shift_wire678),
    .c(shift_wire339)
  );

  wire [5-1:0] shift_wire340;

  muxaltb
  muxcmp340
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire679),
    .b(shift_wire680),
    .c(shift_wire340)
  );

  wire [5-1:0] shift_wire341;

  muxaltb
  muxcmp341
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire681),
    .b(shift_wire682),
    .c(shift_wire341)
  );

  wire [5-1:0] shift_wire342;

  muxaltb
  muxcmp342
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire683),
    .b(shift_wire684),
    .c(shift_wire342)
  );

  wire [5-1:0] shift_wire343;

  muxaltb
  muxcmp343
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire685),
    .b(shift_wire686),
    .c(shift_wire343)
  );

  wire [5-1:0] shift_wire344;

  muxaltb
  muxcmp344
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire687),
    .b(shift_wire688),
    .c(shift_wire344)
  );

  wire [5-1:0] shift_wire345;

  muxaltb
  muxcmp345
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire689),
    .b(shift_wire690),
    .c(shift_wire345)
  );

  wire [5-1:0] shift_wire346;

  muxaltb
  muxcmp346
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire691),
    .b(shift_wire692),
    .c(shift_wire346)
  );

  wire [5-1:0] shift_wire347;

  muxaltb
  muxcmp347
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire693),
    .b(shift_wire694),
    .c(shift_wire347)
  );

  wire [5-1:0] shift_wire348;

  muxaltb
  muxcmp348
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire695),
    .b(shift_wire696),
    .c(shift_wire348)
  );

  wire [5-1:0] shift_wire349;

  muxaltb
  muxcmp349
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire697),
    .b(shift_wire698),
    .c(shift_wire349)
  );

  wire [5-1:0] shift_wire350;

  muxaltb
  muxcmp350
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire699),
    .b(shift_wire700),
    .c(shift_wire350)
  );

  wire [5-1:0] shift_wire351;

  muxaltb
  muxcmp351
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire701),
    .b(shift_wire702),
    .c(shift_wire351)
  );

  wire [5-1:0] shift_wire352;

  muxaltb
  muxcmp352
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire703),
    .b(shift_wire704),
    .c(shift_wire352)
  );

  wire [5-1:0] shift_wire161;

  muxaltb
  muxcmp161
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire321),
    .b(shift_wire322),
    .c(shift_wire161)
  );

  wire [5-1:0] shift_wire162;

  muxaltb
  muxcmp162
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire323),
    .b(shift_wire324),
    .c(shift_wire162)
  );

  wire [5-1:0] shift_wire163;

  muxaltb
  muxcmp163
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire325),
    .b(shift_wire326),
    .c(shift_wire163)
  );

  wire [5-1:0] shift_wire164;

  muxaltb
  muxcmp164
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire327),
    .b(shift_wire328),
    .c(shift_wire164)
  );

  wire [5-1:0] shift_wire165;

  muxaltb
  muxcmp165
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire329),
    .b(shift_wire330),
    .c(shift_wire165)
  );

  wire [5-1:0] shift_wire166;

  muxaltb
  muxcmp166
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire331),
    .b(shift_wire332),
    .c(shift_wire166)
  );

  wire [5-1:0] shift_wire167;

  muxaltb
  muxcmp167
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire333),
    .b(shift_wire334),
    .c(shift_wire167)
  );

  wire [5-1:0] shift_wire168;

  muxaltb
  muxcmp168
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire335),
    .b(shift_wire336),
    .c(shift_wire168)
  );

  wire [5-1:0] shift_wire169;

  muxaltb
  muxcmp169
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire337),
    .b(shift_wire338),
    .c(shift_wire169)
  );

  wire [5-1:0] shift_wire170;

  muxaltb
  muxcmp170
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire339),
    .b(shift_wire340),
    .c(shift_wire170)
  );

  wire [5-1:0] shift_wire171;

  muxaltb
  muxcmp171
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire341),
    .b(shift_wire342),
    .c(shift_wire171)
  );

  wire [5-1:0] shift_wire172;

  muxaltb
  muxcmp172
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire343),
    .b(shift_wire344),
    .c(shift_wire172)
  );

  wire [5-1:0] shift_wire173;

  muxaltb
  muxcmp173
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire345),
    .b(shift_wire346),
    .c(shift_wire173)
  );

  wire [5-1:0] shift_wire174;

  muxaltb
  muxcmp174
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire347),
    .b(shift_wire348),
    .c(shift_wire174)
  );

  wire [5-1:0] shift_wire175;

  muxaltb
  muxcmp175
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire349),
    .b(shift_wire350),
    .c(shift_wire175)
  );

  wire [5-1:0] shift_wire176;

  muxaltb
  muxcmp176
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire351),
    .b(shift_wire352),
    .c(shift_wire176)
  );

  wire [5-1:0] shift_wire81;

  muxaltb
  muxcmp81
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire161),
    .b(shift_wire162),
    .c(shift_wire81)
  );

  wire [5-1:0] shift_wire82;

  muxaltb
  muxcmp82
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire163),
    .b(shift_wire164),
    .c(shift_wire82)
  );

  wire [5-1:0] shift_wire83;

  muxaltb
  muxcmp83
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire165),
    .b(shift_wire166),
    .c(shift_wire83)
  );

  wire [5-1:0] shift_wire84;

  muxaltb
  muxcmp84
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire167),
    .b(shift_wire168),
    .c(shift_wire84)
  );

  wire [5-1:0] shift_wire85;

  muxaltb
  muxcmp85
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire169),
    .b(shift_wire170),
    .c(shift_wire85)
  );

  wire [5-1:0] shift_wire86;

  muxaltb
  muxcmp86
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire171),
    .b(shift_wire172),
    .c(shift_wire86)
  );

  wire [5-1:0] shift_wire87;

  muxaltb
  muxcmp87
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire173),
    .b(shift_wire174),
    .c(shift_wire87)
  );

  wire [5-1:0] shift_wire88;

  muxaltb
  muxcmp88
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire175),
    .b(shift_wire176),
    .c(shift_wire88)
  );

  wire [5-1:0] shift_wire41;

  muxaltb
  muxcmp41
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire81),
    .b(shift_wire82),
    .c(shift_wire41)
  );

  wire [5-1:0] shift_wire42;

  muxaltb
  muxcmp42
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire83),
    .b(shift_wire84),
    .c(shift_wire42)
  );

  wire [5-1:0] shift_wire43;

  muxaltb
  muxcmp43
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire85),
    .b(shift_wire86),
    .c(shift_wire43)
  );

  wire [5-1:0] shift_wire44;

  muxaltb
  muxcmp44
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire87),
    .b(shift_wire88),
    .c(shift_wire44)
  );

  wire [5-1:0] shift_wire21;

  muxaltb
  muxcmp21
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire41),
    .b(shift_wire42),
    .c(shift_wire21)
  );

  wire [5-1:0] shift_wire22;

  muxaltb
  muxcmp22
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire43),
    .b(shift_wire44),
    .c(shift_wire22)
  );

  wire [5-1:0] shift_wire11;

  muxaltb
  muxcmp11
  (
    .clk(clk),
    .rst(rst),
    .a(shift_wire21),
    .b(shift_wire22),
    .c(shift_wire11)
  );

  assign shift_wire = shift_wire11;

endmodule



module muxaltb
(
  input clk,
  input rst,
  input [5-1:0] a,
  input [5-1:0] b,
  output reg [5-1:0] c
);


  always @(posedge clk) begin
    if(rst) begin
      c <= 0;
    end else begin
      if(a < b) begin
        c <= a;
      end else begin
        c <= b;
      end
    end
  end


endmodule

