

module NFA
(
  input clk,
  input rst,
  input [312-1:0] datain,
  output reg [11-1:0] dout
);

  wire [32-1:0] comp;
  wire [76-1:0] w0;
  assign w0[0] = |(datain[311:308] ^ 2);
  assign w0[1] = |(datain[307:304] ^ 1);
  assign w0[2] = |(datain[303:300] ^ 11);
  assign w0[3] = |(datain[299:296] ^ 8);
  assign w0[4] = |(datain[295:292] ^ 0);
  assign w0[5] = |(datain[291:288] ^ 0);
  assign w0[6] = |(datain[287:284] ^ 4);
  assign w0[7] = |(datain[283:280] ^ 2);
  assign w0[8] = |(datain[279:276] ^ 3);
  assign w0[9] = |(datain[275:272] ^ 3);
  assign w0[10] = |(datain[271:268] ^ 12);
  assign w0[11] = |(datain[267:264] ^ 9);
  assign w0[12] = |(datain[263:260] ^ 9);
  assign w0[13] = |(datain[259:256] ^ 9);
  assign w0[14] = |(datain[255:252] ^ 12);
  assign w0[15] = |(datain[251:248] ^ 13);
  assign w0[16] = |(datain[247:244] ^ 2);
  assign w0[17] = |(datain[243:240] ^ 1);
  assign w0[18] = |(datain[239:236] ^ 8);
  assign w0[19] = |(datain[235:232] ^ 11);
  assign w0[20] = |(datain[231:228] ^ 13);
  assign w0[21] = |(datain[227:224] ^ 6);
  assign w0[22] = |(datain[223:220] ^ 11);
  assign w0[23] = |(datain[219:216] ^ 9);
  assign w0[24] = |(datain[215:212] ^ 0);
  assign w0[25] = |(datain[211:208] ^ 3);
  assign w0[26] = |(datain[207:204] ^ 0);
  assign w0[27] = |(datain[203:200] ^ 0);
  assign w0[28] = |(datain[199:196] ^ 11);
  assign w0[29] = |(datain[195:192] ^ 4);
  assign w0[30] = |(datain[191:188] ^ 4);
  assign w0[31] = |(datain[187:184] ^ 0);
  assign w0[32] = |(datain[183:180] ^ 12);
  assign w0[33] = |(datain[179:176] ^ 13);
  assign w0[34] = |(datain[175:172] ^ 2);
  assign w0[35] = |(datain[171:168] ^ 1);
  assign w0[36] = |(datain[167:164] ^ 8);
  assign w0[37] = |(datain[163:160] ^ 11);
  assign w0[38] = |(datain[159:156] ^ 4);
  assign w0[39] = |(datain[155:152] ^ 12);
  assign w0[40] = |(datain[151:148] ^ 1);
  assign w0[41] = |(datain[147:144] ^ 9);
  assign w0[42] = |(datain[143:140] ^ 8);
  assign w0[43] = |(datain[139:136] ^ 11);
  assign w0[44] = |(datain[135:132] ^ 5);
  assign w0[45] = |(datain[131:128] ^ 4);
  assign w0[46] = |(datain[127:124] ^ 1);
  assign w0[47] = |(datain[123:120] ^ 11);
  assign w0[48] = |(datain[119:116] ^ 11);
  assign w0[49] = |(datain[115:112] ^ 8);
  assign w0[50] = |(datain[111:108] ^ 0);
  assign w0[51] = |(datain[107:104] ^ 1);
  assign w0[52] = |(datain[103:100] ^ 5);
  assign w0[53] = |(datain[99:96] ^ 7);
  assign w0[54] = |(datain[95:92] ^ 12);
  assign w0[55] = |(datain[91:88] ^ 13);
  assign w0[56] = |(datain[87:84] ^ 2);
  assign w0[57] = |(datain[83:80] ^ 1);
  assign w0[58] = |(datain[79:76] ^ 11);
  assign w0[59] = |(datain[75:72] ^ 4);
  assign w0[60] = |(datain[71:68] ^ 3);
  assign w0[61] = |(datain[67:64] ^ 14);
  assign w0[62] = |(datain[63:60] ^ 12);
  assign w0[63] = |(datain[59:56] ^ 13);
  assign w0[64] = |(datain[55:52] ^ 2);
  assign w0[65] = |(datain[51:48] ^ 1);
  assign w0[66] = |(datain[47:44] ^ 3);
  assign w0[67] = |(datain[43:40] ^ 2);
  assign w0[68] = |(datain[39:36] ^ 14);
  assign w0[69] = |(datain[35:32] ^ 13);
  assign w0[70] = |(datain[31:28] ^ 8);
  assign w0[71] = |(datain[27:24] ^ 10);
  assign w0[72] = |(datain[23:20] ^ 4);
  assign w0[73] = |(datain[19:16] ^ 12);
  assign w0[74] = |(datain[15:12] ^ 1);
  assign w0[75] = |(datain[11:8] ^ 8);
  assign comp[0] = ~(|w0);
  wire [74-1:0] w1;
  assign w1[0] = |(datain[311:308] ^ 14);
  assign w1[1] = |(datain[307:304] ^ 14);
  assign w1[2] = |(datain[303:300] ^ 5);
  assign w1[3] = |(datain[299:296] ^ 0);
  assign w1[4] = |(datain[295:292] ^ 15);
  assign w1[5] = |(datain[291:288] ^ 7);
  assign w1[6] = |(datain[287:284] ^ 13);
  assign w1[7] = |(datain[283:280] ^ 8);
  assign w1[8] = |(datain[279:276] ^ 2);
  assign w1[9] = |(datain[275:272] ^ 5);
  assign w1[10] = |(datain[271:268] ^ 0);
  assign w1[11] = |(datain[267:264] ^ 15);
  assign w1[12] = |(datain[263:260] ^ 0);
  assign w1[13] = |(datain[259:256] ^ 0);
  assign w1[14] = |(datain[255:252] ^ 8);
  assign w1[15] = |(datain[251:248] ^ 11);
  assign w1[16] = |(datain[247:244] ^ 12);
  assign w1[17] = |(datain[243:240] ^ 8);
  assign w1[18] = |(datain[239:236] ^ 5);
  assign w1[19] = |(datain[235:232] ^ 8);
  assign w1[20] = |(datain[231:228] ^ 0);
  assign w1[21] = |(datain[227:224] ^ 3);
  assign w1[22] = |(datain[223:220] ^ 12);
  assign w1[23] = |(datain[219:216] ^ 1);
  assign w1[24] = |(datain[215:212] ^ 5);
  assign w1[25] = |(datain[211:208] ^ 0);
  assign w1[26] = |(datain[207:204] ^ 11);
  assign w1[27] = |(datain[203:200] ^ 4);
  assign w1[28] = |(datain[199:196] ^ 4);
  assign w1[29] = |(datain[195:192] ^ 0);
  assign w1[30] = |(datain[191:188] ^ 12);
  assign w1[31] = |(datain[187:184] ^ 13);
  assign w1[32] = |(datain[183:180] ^ 2);
  assign w1[33] = |(datain[179:176] ^ 1);
  assign w1[34] = |(datain[175:172] ^ 5);
  assign w1[35] = |(datain[171:168] ^ 8);
  assign w1[36] = |(datain[167:164] ^ 2);
  assign w1[37] = |(datain[163:160] ^ 13);
  assign w1[38] = |(datain[159:156] ^ 0);
  assign w1[39] = |(datain[155:152] ^ 3);
  assign w1[40] = |(datain[151:148] ^ 0);
  assign w1[41] = |(datain[147:144] ^ 0);
  assign w1[42] = |(datain[143:140] ^ 12);
  assign w1[43] = |(datain[139:136] ^ 6);
  assign w1[44] = |(datain[135:132] ^ 0);
  assign w1[45] = |(datain[131:128] ^ 4);
  assign w1[46] = |(datain[127:124] ^ 14);
  assign w1[47] = |(datain[123:120] ^ 9);
  assign w1[48] = |(datain[119:116] ^ 8);
  assign w1[49] = |(datain[115:112] ^ 9);
  assign w1[50] = |(datain[111:108] ^ 4);
  assign w1[51] = |(datain[107:104] ^ 4);
  assign w1[52] = |(datain[103:100] ^ 0);
  assign w1[53] = |(datain[99:96] ^ 1);
  assign w1[54] = |(datain[95:92] ^ 8);
  assign w1[55] = |(datain[91:88] ^ 11);
  assign w1[56] = |(datain[87:84] ^ 13);
  assign w1[57] = |(datain[83:80] ^ 6);
  assign w1[58] = |(datain[79:76] ^ 11);
  assign w1[59] = |(datain[75:72] ^ 9);
  assign w1[60] = |(datain[71:68] ^ 8);
  assign w1[61] = |(datain[67:64] ^ 5);
  assign w1[62] = |(datain[63:60] ^ 0);
  assign w1[63] = |(datain[59:56] ^ 9);
  assign w1[64] = |(datain[55:52] ^ 2);
  assign w1[65] = |(datain[51:48] ^ 11);
  assign w1[66] = |(datain[47:44] ^ 13);
  assign w1[67] = |(datain[43:40] ^ 1);
  assign w1[68] = |(datain[39:36] ^ 0);
  assign w1[69] = |(datain[35:32] ^ 5);
  assign w1[70] = |(datain[31:28] ^ 0);
  assign w1[71] = |(datain[27:24] ^ 3);
  assign w1[72] = |(datain[23:20] ^ 0);
  assign w1[73] = |(datain[19:16] ^ 1);
  assign comp[1] = ~(|w1);
  wire [74-1:0] w2;
  assign w2[0] = |(datain[311:308] ^ 8);
  assign w2[1] = |(datain[307:304] ^ 11);
  assign w2[2] = |(datain[303:300] ^ 14);
  assign w2[3] = |(datain[299:296] ^ 12);
  assign w2[4] = |(datain[295:292] ^ 12);
  assign w2[5] = |(datain[291:288] ^ 7);
  assign w2[6] = |(datain[287:284] ^ 4);
  assign w2[7] = |(datain[283:280] ^ 6);
  assign w2[8] = |(datain[279:276] ^ 0);
  assign w2[9] = |(datain[275:272] ^ 2);
  assign w2[10] = |(datain[271:268] ^ 0);
  assign w2[11] = |(datain[267:264] ^ 0);
  assign w2[12] = |(datain[263:260] ^ 4);
  assign w2[13] = |(datain[259:256] ^ 0);
  assign w2[14] = |(datain[255:252] ^ 5);
  assign w2[15] = |(datain[251:248] ^ 13);
  assign w2[16] = |(datain[247:244] ^ 5);
  assign w2[17] = |(datain[243:240] ^ 8);
  assign w2[18] = |(datain[239:236] ^ 11);
  assign w2[19] = |(datain[235:232] ^ 9);
  assign w2[20] = |(datain[231:228] ^ 0);
  assign w2[21] = |(datain[227:224] ^ 4);
  assign w2[22] = |(datain[223:220] ^ 0);
  assign w2[23] = |(datain[219:216] ^ 0);
  assign w2[24] = |(datain[215:212] ^ 11);
  assign w2[25] = |(datain[211:208] ^ 10);
  assign w2[26] = |(datain[207:204] ^ 4);
  assign w2[27] = |(datain[203:200] ^ 10);
  assign w2[28] = |(datain[199:196] ^ 0);
  assign w2[29] = |(datain[195:192] ^ 8);
  assign w2[30] = |(datain[191:188] ^ 12);
  assign w2[31] = |(datain[187:184] ^ 13);
  assign w2[32] = |(datain[183:180] ^ 2);
  assign w2[33] = |(datain[179:176] ^ 1);
  assign w2[34] = |(datain[175:172] ^ 14);
  assign w2[35] = |(datain[171:168] ^ 9);
  assign w2[36] = |(datain[167:164] ^ 0);
  assign w2[37] = |(datain[163:160] ^ 0);
  assign w2[38] = |(datain[159:156] ^ 0);
  assign w2[39] = |(datain[155:152] ^ 1);
  assign w2[40] = |(datain[151:148] ^ 8);
  assign w2[41] = |(datain[147:144] ^ 0);
  assign w2[42] = |(datain[143:140] ^ 3);
  assign w2[43] = |(datain[139:136] ^ 14);
  assign w2[44] = |(datain[135:132] ^ 6);
  assign w2[45] = |(datain[131:128] ^ 2);
  assign w2[46] = |(datain[127:124] ^ 0);
  assign w2[47] = |(datain[123:120] ^ 8);
  assign w2[48] = |(datain[119:116] ^ 4);
  assign w2[49] = |(datain[115:112] ^ 0);
  assign w2[50] = |(datain[111:108] ^ 7);
  assign w2[51] = |(datain[107:104] ^ 4);
  assign w2[52] = |(datain[103:100] ^ 1);
  assign w2[53] = |(datain[99:96] ^ 1);
  assign w2[54] = |(datain[95:92] ^ 8);
  assign w2[55] = |(datain[91:88] ^ 0);
  assign w2[56] = |(datain[87:84] ^ 3);
  assign w2[57] = |(datain[83:80] ^ 14);
  assign w2[58] = |(datain[79:76] ^ 5);
  assign w2[59] = |(datain[75:72] ^ 12);
  assign w2[60] = |(datain[71:68] ^ 0);
  assign w2[61] = |(datain[67:64] ^ 8);
  assign w2[62] = |(datain[63:60] ^ 6);
  assign w2[63] = |(datain[59:56] ^ 11);
  assign w2[64] = |(datain[55:52] ^ 7);
  assign w2[65] = |(datain[51:48] ^ 4);
  assign w2[66] = |(datain[47:44] ^ 0);
  assign w2[67] = |(datain[43:40] ^ 10);
  assign w2[68] = |(datain[39:36] ^ 10);
  assign w2[69] = |(datain[35:32] ^ 1);
  assign w2[70] = |(datain[31:28] ^ 4);
  assign w2[71] = |(datain[27:24] ^ 10);
  assign w2[72] = |(datain[23:20] ^ 0);
  assign w2[73] = |(datain[19:16] ^ 8);
  assign comp[2] = ~(|w2);
  wire [74-1:0] w3;
  assign w3[0] = |(datain[311:308] ^ 5);
  assign w3[1] = |(datain[307:304] ^ 5);
  assign w3[2] = |(datain[303:300] ^ 8);
  assign w3[3] = |(datain[299:296] ^ 11);
  assign w3[4] = |(datain[295:292] ^ 14);
  assign w3[5] = |(datain[291:288] ^ 12);
  assign w3[6] = |(datain[287:284] ^ 12);
  assign w3[7] = |(datain[283:280] ^ 7);
  assign w3[8] = |(datain[279:276] ^ 4);
  assign w3[9] = |(datain[275:272] ^ 6);
  assign w3[10] = |(datain[271:268] ^ 0);
  assign w3[11] = |(datain[267:264] ^ 2);
  assign w3[12] = |(datain[263:260] ^ 0);
  assign w3[13] = |(datain[259:256] ^ 0);
  assign w3[14] = |(datain[255:252] ^ 4);
  assign w3[15] = |(datain[251:248] ^ 0);
  assign w3[16] = |(datain[247:244] ^ 5);
  assign w3[17] = |(datain[243:240] ^ 13);
  assign w3[18] = |(datain[239:236] ^ 5);
  assign w3[19] = |(datain[235:232] ^ 8);
  assign w3[20] = |(datain[231:228] ^ 3);
  assign w3[21] = |(datain[227:224] ^ 3);
  assign w3[22] = |(datain[223:220] ^ 13);
  assign w3[23] = |(datain[219:216] ^ 2);
  assign w3[24] = |(datain[215:212] ^ 11);
  assign w3[25] = |(datain[211:208] ^ 9);
  assign w3[26] = |(datain[207:204] ^ 8);
  assign w3[27] = |(datain[203:200] ^ 7);
  assign w3[28] = |(datain[199:196] ^ 0);
  assign w3[29] = |(datain[195:192] ^ 0);
  assign w3[30] = |(datain[191:188] ^ 12);
  assign w3[31] = |(datain[187:184] ^ 13);
  assign w3[32] = |(datain[183:180] ^ 2);
  assign w3[33] = |(datain[179:176] ^ 1);
  assign w3[34] = |(datain[175:172] ^ 5);
  assign w3[35] = |(datain[171:168] ^ 0);
  assign w3[36] = |(datain[167:164] ^ 5);
  assign w3[37] = |(datain[163:160] ^ 5);
  assign w3[38] = |(datain[159:156] ^ 8);
  assign w3[39] = |(datain[155:152] ^ 11);
  assign w3[40] = |(datain[151:148] ^ 14);
  assign w3[41] = |(datain[147:144] ^ 12);
  assign w3[42] = |(datain[143:140] ^ 12);
  assign w3[43] = |(datain[139:136] ^ 7);
  assign w3[44] = |(datain[135:132] ^ 4);
  assign w3[45] = |(datain[131:128] ^ 6);
  assign w3[46] = |(datain[127:124] ^ 0);
  assign w3[47] = |(datain[123:120] ^ 2);
  assign w3[48] = |(datain[119:116] ^ 0);
  assign w3[49] = |(datain[115:112] ^ 0);
  assign w3[50] = |(datain[111:108] ^ 4);
  assign w3[51] = |(datain[107:104] ^ 0);
  assign w3[52] = |(datain[103:100] ^ 5);
  assign w3[53] = |(datain[99:96] ^ 13);
  assign w3[54] = |(datain[95:92] ^ 5);
  assign w3[55] = |(datain[91:88] ^ 8);
  assign w3[56] = |(datain[87:84] ^ 11);
  assign w3[57] = |(datain[83:80] ^ 10);
  assign w3[58] = |(datain[79:76] ^ 9);
  assign w3[59] = |(datain[75:72] ^ 10);
  assign w3[60] = |(datain[71:68] ^ 1);
  assign w3[61] = |(datain[67:64] ^ 0);
  assign w3[62] = |(datain[63:60] ^ 11);
  assign w3[63] = |(datain[59:56] ^ 9);
  assign w3[64] = |(datain[55:52] ^ 1);
  assign w3[65] = |(datain[51:48] ^ 3);
  assign w3[66] = |(datain[47:44] ^ 1);
  assign w3[67] = |(datain[43:40] ^ 0);
  assign w3[68] = |(datain[39:36] ^ 12);
  assign w3[69] = |(datain[35:32] ^ 13);
  assign w3[70] = |(datain[31:28] ^ 2);
  assign w3[71] = |(datain[27:24] ^ 1);
  assign w3[72] = |(datain[23:20] ^ 11);
  assign w3[73] = |(datain[19:16] ^ 8);
  assign comp[3] = ~(|w3);
  wire [74-1:0] w4;
  assign w4[0] = |(datain[311:308] ^ 8);
  assign w4[1] = |(datain[307:304] ^ 11);
  assign w4[2] = |(datain[303:300] ^ 14);
  assign w4[3] = |(datain[299:296] ^ 12);
  assign w4[4] = |(datain[295:292] ^ 12);
  assign w4[5] = |(datain[291:288] ^ 7);
  assign w4[6] = |(datain[287:284] ^ 4);
  assign w4[7] = |(datain[283:280] ^ 6);
  assign w4[8] = |(datain[279:276] ^ 0);
  assign w4[9] = |(datain[275:272] ^ 2);
  assign w4[10] = |(datain[271:268] ^ 0);
  assign w4[11] = |(datain[267:264] ^ 0);
  assign w4[12] = |(datain[263:260] ^ 4);
  assign w4[13] = |(datain[259:256] ^ 0);
  assign w4[14] = |(datain[255:252] ^ 5);
  assign w4[15] = |(datain[251:248] ^ 13);
  assign w4[16] = |(datain[247:244] ^ 5);
  assign w4[17] = |(datain[243:240] ^ 8);
  assign w4[18] = |(datain[239:236] ^ 11);
  assign w4[19] = |(datain[235:232] ^ 10);
  assign w4[20] = |(datain[231:228] ^ 9);
  assign w4[21] = |(datain[227:224] ^ 10);
  assign w4[22] = |(datain[223:220] ^ 1);
  assign w4[23] = |(datain[219:216] ^ 0);
  assign w4[24] = |(datain[215:212] ^ 11);
  assign w4[25] = |(datain[211:208] ^ 9);
  assign w4[26] = |(datain[207:204] ^ 1);
  assign w4[27] = |(datain[203:200] ^ 3);
  assign w4[28] = |(datain[199:196] ^ 1);
  assign w4[29] = |(datain[195:192] ^ 0);
  assign w4[30] = |(datain[191:188] ^ 12);
  assign w4[31] = |(datain[187:184] ^ 13);
  assign w4[32] = |(datain[183:180] ^ 2);
  assign w4[33] = |(datain[179:176] ^ 1);
  assign w4[34] = |(datain[175:172] ^ 11);
  assign w4[35] = |(datain[171:168] ^ 8);
  assign w4[36] = |(datain[167:164] ^ 0);
  assign w4[37] = |(datain[163:160] ^ 0);
  assign w4[38] = |(datain[159:156] ^ 4);
  assign w4[39] = |(datain[155:152] ^ 2);
  assign w4[40] = |(datain[151:148] ^ 5);
  assign w4[41] = |(datain[147:144] ^ 0);
  assign w4[42] = |(datain[143:140] ^ 5);
  assign w4[43] = |(datain[139:136] ^ 8);
  assign w4[44] = |(datain[135:132] ^ 3);
  assign w4[45] = |(datain[131:128] ^ 3);
  assign w4[46] = |(datain[127:124] ^ 12);
  assign w4[47] = |(datain[123:120] ^ 9);
  assign w4[48] = |(datain[119:116] ^ 3);
  assign w4[49] = |(datain[115:112] ^ 3);
  assign w4[50] = |(datain[111:108] ^ 13);
  assign w4[51] = |(datain[107:104] ^ 2);
  assign w4[52] = |(datain[103:100] ^ 12);
  assign w4[53] = |(datain[99:96] ^ 13);
  assign w4[54] = |(datain[95:92] ^ 2);
  assign w4[55] = |(datain[91:88] ^ 1);
  assign w4[56] = |(datain[87:84] ^ 5);
  assign w4[57] = |(datain[83:80] ^ 0);
  assign w4[58] = |(datain[79:76] ^ 5);
  assign w4[59] = |(datain[75:72] ^ 5);
  assign w4[60] = |(datain[71:68] ^ 8);
  assign w4[61] = |(datain[67:64] ^ 11);
  assign w4[62] = |(datain[63:60] ^ 14);
  assign w4[63] = |(datain[59:56] ^ 12);
  assign w4[64] = |(datain[55:52] ^ 12);
  assign w4[65] = |(datain[51:48] ^ 7);
  assign w4[66] = |(datain[47:44] ^ 4);
  assign w4[67] = |(datain[43:40] ^ 6);
  assign w4[68] = |(datain[39:36] ^ 0);
  assign w4[69] = |(datain[35:32] ^ 2);
  assign w4[70] = |(datain[31:28] ^ 0);
  assign w4[71] = |(datain[27:24] ^ 0);
  assign w4[72] = |(datain[23:20] ^ 4);
  assign w4[73] = |(datain[19:16] ^ 0);
  assign comp[4] = ~(|w4);
  wire [76-1:0] w5;
  assign w5[0] = |(datain[311:308] ^ 12);
  assign w5[1] = |(datain[307:304] ^ 13);
  assign w5[2] = |(datain[303:300] ^ 2);
  assign w5[3] = |(datain[299:296] ^ 1);
  assign w5[4] = |(datain[295:292] ^ 3);
  assign w5[5] = |(datain[291:288] ^ 3);
  assign w5[6] = |(datain[287:284] ^ 12);
  assign w5[7] = |(datain[283:280] ^ 9);
  assign w5[8] = |(datain[279:276] ^ 11);
  assign w5[9] = |(datain[275:272] ^ 8);
  assign w5[10] = |(datain[271:268] ^ 0);
  assign w5[11] = |(datain[267:264] ^ 0);
  assign w5[12] = |(datain[263:260] ^ 4);
  assign w5[13] = |(datain[259:256] ^ 2);
  assign w5[14] = |(datain[255:252] ^ 9);
  assign w5[15] = |(datain[251:248] ^ 9);
  assign w5[16] = |(datain[247:244] ^ 12);
  assign w5[17] = |(datain[243:240] ^ 13);
  assign w5[18] = |(datain[239:236] ^ 2);
  assign w5[19] = |(datain[235:232] ^ 1);
  assign w5[20] = |(datain[231:228] ^ 11);
  assign w5[21] = |(datain[227:224] ^ 4);
  assign w5[22] = |(datain[223:220] ^ 4);
  assign w5[23] = |(datain[219:216] ^ 0);
  assign w5[24] = |(datain[215:212] ^ 11);
  assign w5[25] = |(datain[211:208] ^ 10);
  assign w5[26] = |(datain[207:204] ^ 8);
  assign w5[27] = |(datain[203:200] ^ 9);
  assign w5[28] = |(datain[199:196] ^ 0);
  assign w5[29] = |(datain[195:192] ^ 4);
  assign w5[30] = |(datain[191:188] ^ 5);
  assign w5[31] = |(datain[187:184] ^ 9);
  assign w5[32] = |(datain[183:180] ^ 12);
  assign w5[33] = |(datain[179:176] ^ 13);
  assign w5[34] = |(datain[175:172] ^ 2);
  assign w5[35] = |(datain[171:168] ^ 1);
  assign w5[36] = |(datain[167:164] ^ 11);
  assign w5[37] = |(datain[163:160] ^ 8);
  assign w5[38] = |(datain[159:156] ^ 0);
  assign w5[39] = |(datain[155:152] ^ 1);
  assign w5[40] = |(datain[151:148] ^ 5);
  assign w5[41] = |(datain[147:144] ^ 7);
  assign w5[42] = |(datain[143:140] ^ 5);
  assign w5[43] = |(datain[139:136] ^ 10);
  assign w5[44] = |(datain[135:132] ^ 5);
  assign w5[45] = |(datain[131:128] ^ 9);
  assign w5[46] = |(datain[127:124] ^ 12);
  assign w5[47] = |(datain[123:120] ^ 13);
  assign w5[48] = |(datain[119:116] ^ 2);
  assign w5[49] = |(datain[115:112] ^ 1);
  assign w5[50] = |(datain[111:108] ^ 11);
  assign w5[51] = |(datain[107:104] ^ 4);
  assign w5[52] = |(datain[103:100] ^ 3);
  assign w5[53] = |(datain[99:96] ^ 14);
  assign w5[54] = |(datain[95:92] ^ 12);
  assign w5[55] = |(datain[91:88] ^ 13);
  assign w5[56] = |(datain[87:84] ^ 2);
  assign w5[57] = |(datain[83:80] ^ 1);
  assign w5[58] = |(datain[79:76] ^ 5);
  assign w5[59] = |(datain[75:72] ^ 8);
  assign w5[60] = |(datain[71:68] ^ 5);
  assign w5[61] = |(datain[67:64] ^ 10);
  assign w5[62] = |(datain[63:60] ^ 1);
  assign w5[63] = |(datain[59:56] ^ 15);
  assign w5[64] = |(datain[55:52] ^ 5);
  assign w5[65] = |(datain[51:48] ^ 9);
  assign w5[66] = |(datain[47:44] ^ 12);
  assign w5[67] = |(datain[43:40] ^ 13);
  assign w5[68] = |(datain[39:36] ^ 2);
  assign w5[69] = |(datain[35:32] ^ 1);
  assign w5[70] = |(datain[31:28] ^ 5);
  assign w5[71] = |(datain[27:24] ^ 10);
  assign w5[72] = |(datain[23:20] ^ 1);
  assign w5[73] = |(datain[19:16] ^ 15);
  assign w5[74] = |(datain[15:12] ^ 11);
  assign w5[75] = |(datain[11:8] ^ 8);
  assign comp[5] = ~(|w5);
  wire [76-1:0] w6;
  assign w6[0] = |(datain[311:308] ^ 8);
  assign w6[1] = |(datain[307:304] ^ 9);
  assign w6[2] = |(datain[303:300] ^ 4);
  assign w6[3] = |(datain[299:296] ^ 5);
  assign w6[4] = |(datain[295:292] ^ 1);
  assign w6[5] = |(datain[291:288] ^ 5);
  assign w6[6] = |(datain[287:284] ^ 5);
  assign w6[7] = |(datain[283:280] ^ 0);
  assign w6[8] = |(datain[279:276] ^ 5);
  assign w6[9] = |(datain[275:272] ^ 6);
  assign w6[10] = |(datain[271:268] ^ 5);
  assign w6[11] = |(datain[267:264] ^ 7);
  assign w6[12] = |(datain[263:260] ^ 5);
  assign w6[13] = |(datain[259:256] ^ 5);
  assign w6[14] = |(datain[255:252] ^ 1);
  assign w6[15] = |(datain[251:248] ^ 14);
  assign w6[16] = |(datain[247:244] ^ 0);
  assign w6[17] = |(datain[243:240] ^ 6);
  assign w6[18] = |(datain[239:236] ^ 5);
  assign w6[19] = |(datain[235:232] ^ 3);
  assign w6[20] = |(datain[231:228] ^ 14);
  assign w6[21] = |(datain[227:224] ^ 8);
  assign w6[22] = |(datain[223:220] ^ 4);
  assign w6[23] = |(datain[219:216] ^ 12);
  assign w6[24] = |(datain[215:212] ^ 0);
  assign w6[25] = |(datain[211:208] ^ 0);
  assign w6[26] = |(datain[207:204] ^ 5);
  assign w6[27] = |(datain[203:200] ^ 11);
  assign w6[28] = |(datain[199:196] ^ 11);
  assign w6[29] = |(datain[195:192] ^ 4);
  assign w6[30] = |(datain[191:188] ^ 4);
  assign w6[31] = |(datain[187:184] ^ 0);
  assign w6[32] = |(datain[183:180] ^ 12);
  assign w6[33] = |(datain[179:176] ^ 13);
  assign w6[34] = |(datain[175:172] ^ 2);
  assign w6[35] = |(datain[171:168] ^ 1);
  assign w6[36] = |(datain[167:164] ^ 3);
  assign w6[37] = |(datain[163:160] ^ 11);
  assign w6[38] = |(datain[159:156] ^ 12);
  assign w6[39] = |(datain[155:152] ^ 8);
  assign w6[40] = |(datain[151:148] ^ 0);
  assign w6[41] = |(datain[147:144] ^ 7);
  assign w6[42] = |(datain[143:140] ^ 1);
  assign w6[43] = |(datain[139:136] ^ 15);
  assign w6[44] = |(datain[135:132] ^ 5);
  assign w6[45] = |(datain[131:128] ^ 13);
  assign w6[46] = |(datain[127:124] ^ 5);
  assign w6[47] = |(datain[123:120] ^ 15);
  assign w6[48] = |(datain[119:116] ^ 5);
  assign w6[49] = |(datain[115:112] ^ 14);
  assign w6[50] = |(datain[111:108] ^ 5);
  assign w6[51] = |(datain[107:104] ^ 8);
  assign w6[52] = |(datain[103:100] ^ 7);
  assign w6[53] = |(datain[99:96] ^ 5);
  assign w6[54] = |(datain[95:92] ^ 1);
  assign w6[55] = |(datain[91:88] ^ 9);
  assign w6[56] = |(datain[87:84] ^ 12);
  assign w6[57] = |(datain[83:80] ^ 7);
  assign w6[58] = |(datain[79:76] ^ 0);
  assign w6[59] = |(datain[75:72] ^ 4);
  assign w6[60] = |(datain[71:68] ^ 4);
  assign w6[61] = |(datain[67:64] ^ 13);
  assign w6[62] = |(datain[63:60] ^ 14);
  assign w6[63] = |(datain[59:56] ^ 9);
  assign w6[64] = |(datain[55:52] ^ 2);
  assign w6[65] = |(datain[51:48] ^ 13);
  assign w6[66] = |(datain[47:44] ^ 0);
  assign w6[67] = |(datain[43:40] ^ 4);
  assign w6[68] = |(datain[39:36] ^ 0);
  assign w6[69] = |(datain[35:32] ^ 0);
  assign w6[70] = |(datain[31:28] ^ 8);
  assign w6[71] = |(datain[27:24] ^ 9);
  assign w6[72] = |(datain[23:20] ^ 4);
  assign w6[73] = |(datain[19:16] ^ 4);
  assign w6[74] = |(datain[15:12] ^ 0);
  assign w6[75] = |(datain[11:8] ^ 2);
  assign comp[6] = ~(|w6);
  wire [76-1:0] w7;
  assign w7[0] = |(datain[311:308] ^ 8);
  assign w7[1] = |(datain[307:304] ^ 9);
  assign w7[2] = |(datain[303:300] ^ 4);
  assign w7[3] = |(datain[299:296] ^ 4);
  assign w7[4] = |(datain[295:292] ^ 0);
  assign w7[5] = |(datain[291:288] ^ 2);
  assign w7[6] = |(datain[287:284] ^ 3);
  assign w7[7] = |(datain[283:280] ^ 3);
  assign w7[8] = |(datain[279:276] ^ 12);
  assign w7[9] = |(datain[275:272] ^ 0);
  assign w7[10] = |(datain[271:268] ^ 2);
  assign w7[11] = |(datain[267:264] ^ 6);
  assign w7[12] = |(datain[263:260] ^ 8);
  assign w7[13] = |(datain[259:256] ^ 9);
  assign w7[14] = |(datain[255:252] ^ 4);
  assign w7[15] = |(datain[251:248] ^ 5);
  assign w7[16] = |(datain[247:244] ^ 1);
  assign w7[17] = |(datain[243:240] ^ 5);
  assign w7[18] = |(datain[239:236] ^ 11);
  assign w7[19] = |(datain[235:232] ^ 9);
  assign w7[20] = |(datain[231:228] ^ 0);
  assign w7[21] = |(datain[227:224] ^ 4);
  assign w7[22] = |(datain[223:220] ^ 0);
  assign w7[23] = |(datain[219:216] ^ 0);
  assign w7[24] = |(datain[215:212] ^ 8);
  assign w7[25] = |(datain[211:208] ^ 11);
  assign w7[26] = |(datain[207:204] ^ 13);
  assign w7[27] = |(datain[203:200] ^ 6);
  assign w7[28] = |(datain[199:196] ^ 11);
  assign w7[29] = |(datain[195:192] ^ 4);
  assign w7[30] = |(datain[191:188] ^ 4);
  assign w7[31] = |(datain[187:184] ^ 0);
  assign w7[32] = |(datain[183:180] ^ 12);
  assign w7[33] = |(datain[179:176] ^ 13);
  assign w7[34] = |(datain[175:172] ^ 2);
  assign w7[35] = |(datain[171:168] ^ 1);
  assign w7[36] = |(datain[167:164] ^ 0);
  assign w7[37] = |(datain[163:160] ^ 6);
  assign w7[38] = |(datain[159:156] ^ 1);
  assign w7[39] = |(datain[155:152] ^ 15);
  assign w7[40] = |(datain[151:148] ^ 8);
  assign w7[41] = |(datain[147:144] ^ 15);
  assign w7[42] = |(datain[143:140] ^ 4);
  assign w7[43] = |(datain[139:136] ^ 5);
  assign w7[44] = |(datain[135:132] ^ 1);
  assign w7[45] = |(datain[131:128] ^ 5);
  assign w7[46] = |(datain[127:124] ^ 8);
  assign w7[47] = |(datain[123:120] ^ 0);
  assign w7[48] = |(datain[119:116] ^ 4);
  assign w7[49] = |(datain[115:112] ^ 13);
  assign w7[50] = |(datain[111:108] ^ 0);
  assign w7[51] = |(datain[107:104] ^ 6);
  assign w7[52] = |(datain[103:100] ^ 4);
  assign w7[53] = |(datain[99:96] ^ 0);
  assign w7[54] = |(datain[95:92] ^ 11);
  assign w7[55] = |(datain[91:88] ^ 4);
  assign w7[56] = |(datain[87:84] ^ 3);
  assign w7[57] = |(datain[83:80] ^ 14);
  assign w7[58] = |(datain[79:76] ^ 9);
  assign w7[59] = |(datain[75:72] ^ 12);
  assign w7[60] = |(datain[71:68] ^ 0);
  assign w7[61] = |(datain[67:64] ^ 14);
  assign w7[62] = |(datain[63:60] ^ 14);
  assign w7[63] = |(datain[59:56] ^ 8);
  assign w7[64] = |(datain[55:52] ^ 13);
  assign w7[65] = |(datain[51:48] ^ 8);
  assign w7[66] = |(datain[47:44] ^ 15);
  assign w7[67] = |(datain[43:40] ^ 14);
  assign w7[68] = |(datain[39:36] ^ 8);
  assign w7[69] = |(datain[35:32] ^ 0);
  assign w7[70] = |(datain[31:28] ^ 4);
  assign w7[71] = |(datain[27:24] ^ 13);
  assign w7[72] = |(datain[23:20] ^ 0);
  assign w7[73] = |(datain[19:16] ^ 5);
  assign w7[74] = |(datain[15:12] ^ 4);
  assign w7[75] = |(datain[11:8] ^ 0);
  assign comp[7] = ~(|w7);
  wire [74-1:0] w8;
  assign w8[0] = |(datain[311:308] ^ 11);
  assign w8[1] = |(datain[307:304] ^ 4);
  assign w8[2] = |(datain[303:300] ^ 4);
  assign w8[3] = |(datain[299:296] ^ 0);
  assign w8[4] = |(datain[295:292] ^ 12);
  assign w8[5] = |(datain[291:288] ^ 13);
  assign w8[6] = |(datain[287:284] ^ 2);
  assign w8[7] = |(datain[283:280] ^ 1);
  assign w8[8] = |(datain[279:276] ^ 14);
  assign w8[9] = |(datain[275:272] ^ 8);
  assign w8[10] = |(datain[271:268] ^ 0);
  assign w8[11] = |(datain[267:264] ^ 13);
  assign w8[12] = |(datain[263:260] ^ 0);
  assign w8[13] = |(datain[259:256] ^ 0);
  assign w8[14] = |(datain[255:252] ^ 11);
  assign w8[15] = |(datain[251:248] ^ 9);
  assign w8[16] = |(datain[247:244] ^ 1);
  assign w8[17] = |(datain[243:240] ^ 8);
  assign w8[18] = |(datain[239:236] ^ 0);
  assign w8[19] = |(datain[235:232] ^ 0);
  assign w8[20] = |(datain[231:228] ^ 11);
  assign w8[21] = |(datain[227:224] ^ 10);
  assign w8[22] = |(datain[223:220] ^ 10);
  assign w8[23] = |(datain[219:216] ^ 7);
  assign w8[24] = |(datain[215:212] ^ 0);
  assign w8[25] = |(datain[211:208] ^ 2);
  assign w8[26] = |(datain[207:204] ^ 11);
  assign w8[27] = |(datain[203:200] ^ 4);
  assign w8[28] = |(datain[199:196] ^ 4);
  assign w8[29] = |(datain[195:192] ^ 0);
  assign w8[30] = |(datain[191:188] ^ 12);
  assign w8[31] = |(datain[187:184] ^ 13);
  assign w8[32] = |(datain[183:180] ^ 2);
  assign w8[33] = |(datain[179:176] ^ 1);
  assign w8[34] = |(datain[175:172] ^ 14);
  assign w8[35] = |(datain[171:168] ^ 9);
  assign w8[36] = |(datain[167:164] ^ 5);
  assign w8[37] = |(datain[163:160] ^ 2);
  assign w8[38] = |(datain[159:156] ^ 15);
  assign w8[39] = |(datain[155:152] ^ 15);
  assign w8[40] = |(datain[151:148] ^ 3);
  assign w8[41] = |(datain[147:144] ^ 2);
  assign w8[42] = |(datain[143:140] ^ 12);
  assign w8[43] = |(datain[139:136] ^ 0);
  assign w8[44] = |(datain[135:132] ^ 14);
  assign w8[45] = |(datain[131:128] ^ 11);
  assign w8[46] = |(datain[127:124] ^ 0);
  assign w8[47] = |(datain[123:120] ^ 2);
  assign w8[48] = |(datain[119:116] ^ 11);
  assign w8[49] = |(datain[115:112] ^ 0);
  assign w8[50] = |(datain[111:108] ^ 0);
  assign w8[51] = |(datain[107:104] ^ 2);
  assign w8[52] = |(datain[103:100] ^ 11);
  assign w8[53] = |(datain[99:96] ^ 4);
  assign w8[54] = |(datain[95:92] ^ 4);
  assign w8[55] = |(datain[91:88] ^ 2);
  assign w8[56] = |(datain[87:84] ^ 3);
  assign w8[57] = |(datain[83:80] ^ 3);
  assign w8[58] = |(datain[79:76] ^ 12);
  assign w8[59] = |(datain[75:72] ^ 9);
  assign w8[60] = |(datain[71:68] ^ 3);
  assign w8[61] = |(datain[67:64] ^ 3);
  assign w8[62] = |(datain[63:60] ^ 13);
  assign w8[63] = |(datain[59:56] ^ 2);
  assign w8[64] = |(datain[55:52] ^ 12);
  assign w8[65] = |(datain[51:48] ^ 13);
  assign w8[66] = |(datain[47:44] ^ 2);
  assign w8[67] = |(datain[43:40] ^ 1);
  assign w8[68] = |(datain[39:36] ^ 12);
  assign w8[69] = |(datain[35:32] ^ 3);
  assign w8[70] = |(datain[31:28] ^ 11);
  assign w8[71] = |(datain[27:24] ^ 15);
  assign w8[72] = |(datain[23:20] ^ 0);
  assign w8[73] = |(datain[19:16] ^ 2);
  assign comp[8] = ~(|w8);
  wire [76-1:0] w9;
  assign w9[0] = |(datain[311:308] ^ 12);
  assign w9[1] = |(datain[307:304] ^ 9);
  assign w9[2] = |(datain[303:300] ^ 8);
  assign w9[3] = |(datain[299:296] ^ 11);
  assign w9[4] = |(datain[295:292] ^ 13);
  assign w9[5] = |(datain[291:288] ^ 1);
  assign w9[6] = |(datain[287:284] ^ 11);
  assign w9[7] = |(datain[283:280] ^ 8);
  assign w9[8] = |(datain[279:276] ^ 0);
  assign w9[9] = |(datain[275:272] ^ 2);
  assign w9[10] = |(datain[271:268] ^ 4);
  assign w9[11] = |(datain[267:264] ^ 2);
  assign w9[12] = |(datain[263:260] ^ 2);
  assign w9[13] = |(datain[259:256] ^ 14);
  assign w9[14] = |(datain[255:252] ^ 8);
  assign w9[15] = |(datain[251:248] ^ 11);
  assign w9[16] = |(datain[247:244] ^ 1);
  assign w9[17] = |(datain[243:240] ^ 14);
  assign w9[18] = |(datain[239:236] ^ 3);
  assign w9[19] = |(datain[235:232] ^ 9);
  assign w9[20] = |(datain[231:228] ^ 0);
  assign w9[21] = |(datain[227:224] ^ 15);
  assign w9[22] = |(datain[223:220] ^ 9);
  assign w9[23] = |(datain[219:216] ^ 12);
  assign w9[24] = |(datain[215:212] ^ 15);
  assign w9[25] = |(datain[211:208] ^ 10);
  assign w9[26] = |(datain[207:204] ^ 2);
  assign w9[27] = |(datain[203:200] ^ 14);
  assign w9[28] = |(datain[199:196] ^ 15);
  assign w9[29] = |(datain[195:192] ^ 15);
  assign w9[30] = |(datain[191:188] ^ 1);
  assign w9[31] = |(datain[187:184] ^ 14);
  assign w9[32] = |(datain[183:180] ^ 14);
  assign w9[33] = |(datain[179:176] ^ 8);
  assign w9[34] = |(datain[175:172] ^ 0);
  assign w9[35] = |(datain[171:168] ^ 13);
  assign w9[36] = |(datain[167:164] ^ 12);
  assign w9[37] = |(datain[163:160] ^ 3);
  assign w9[38] = |(datain[159:156] ^ 8);
  assign w9[39] = |(datain[155:152] ^ 11);
  assign w9[40] = |(datain[151:148] ^ 14);
  assign w9[41] = |(datain[147:144] ^ 12);
  assign w9[42] = |(datain[143:140] ^ 11);
  assign w9[43] = |(datain[139:136] ^ 8);
  assign w9[44] = |(datain[135:132] ^ 0);
  assign w9[45] = |(datain[131:128] ^ 0);
  assign w9[46] = |(datain[127:124] ^ 5);
  assign w9[47] = |(datain[123:120] ^ 7);
  assign w9[48] = |(datain[119:116] ^ 14);
  assign w9[49] = |(datain[115:112] ^ 8);
  assign w9[50] = |(datain[111:108] ^ 14);
  assign w9[51] = |(datain[107:104] ^ 11);
  assign w9[52] = |(datain[103:100] ^ 15);
  assign w9[53] = |(datain[99:96] ^ 15);
  assign w9[54] = |(datain[95:92] ^ 11);
  assign w9[55] = |(datain[91:88] ^ 11);
  assign w9[56] = |(datain[87:84] ^ 6);
  assign w9[57] = |(datain[83:80] ^ 3);
  assign w9[58] = |(datain[79:76] ^ 0);
  assign w9[59] = |(datain[75:72] ^ 15);
  assign w9[60] = |(datain[71:68] ^ 8);
  assign w9[61] = |(datain[67:64] ^ 9);
  assign w9[62] = |(datain[63:60] ^ 0);
  assign w9[63] = |(datain[59:56] ^ 15);
  assign w9[64] = |(datain[55:52] ^ 8);
  assign w9[65] = |(datain[51:48] ^ 9);
  assign w9[66] = |(datain[47:44] ^ 5);
  assign w9[67] = |(datain[43:40] ^ 7);
  assign w9[68] = |(datain[39:36] ^ 0);
  assign w9[69] = |(datain[35:32] ^ 2);
  assign w9[70] = |(datain[31:28] ^ 14);
  assign w9[71] = |(datain[27:24] ^ 8);
  assign w9[72] = |(datain[23:20] ^ 12);
  assign w9[73] = |(datain[19:16] ^ 8);
  assign w9[74] = |(datain[15:12] ^ 0);
  assign w9[75] = |(datain[11:8] ^ 2);
  assign comp[9] = ~(|w9);
  wire [74-1:0] w10;
  assign w10[0] = |(datain[311:308] ^ 0);
  assign w10[1] = |(datain[307:304] ^ 10);
  assign w10[2] = |(datain[303:300] ^ 5);
  assign w10[3] = |(datain[299:296] ^ 2);
  assign w10[4] = |(datain[295:292] ^ 5);
  assign w10[5] = |(datain[291:288] ^ 3);
  assign w10[6] = |(datain[287:284] ^ 5);
  assign w10[7] = |(datain[283:280] ^ 6);
  assign w10[8] = |(datain[279:276] ^ 8);
  assign w10[9] = |(datain[275:272] ^ 11);
  assign w10[10] = |(datain[271:268] ^ 13);
  assign w10[11] = |(datain[267:264] ^ 13);
  assign w10[12] = |(datain[263:260] ^ 15);
  assign w10[13] = |(datain[259:256] ^ 14);
  assign w10[14] = |(datain[255:252] ^ 12);
  assign w10[15] = |(datain[251:248] ^ 7);
  assign w10[16] = |(datain[247:244] ^ 14);
  assign w10[17] = |(datain[243:240] ^ 8);
  assign w10[18] = |(datain[239:236] ^ 13);
  assign w10[19] = |(datain[235:232] ^ 4);
  assign w10[20] = |(datain[231:228] ^ 15);
  assign w10[21] = |(datain[227:224] ^ 7);
  assign w10[22] = |(datain[223:220] ^ 11);
  assign w10[23] = |(datain[219:216] ^ 4);
  assign w10[24] = |(datain[215:212] ^ 4);
  assign w10[25] = |(datain[211:208] ^ 0);
  assign w10[26] = |(datain[207:204] ^ 5);
  assign w10[27] = |(datain[203:200] ^ 10);
  assign w10[28] = |(datain[199:196] ^ 5);
  assign w10[29] = |(datain[195:192] ^ 11);
  assign w10[30] = |(datain[191:188] ^ 12);
  assign w10[31] = |(datain[187:184] ^ 13);
  assign w10[32] = |(datain[183:180] ^ 2);
  assign w10[33] = |(datain[179:176] ^ 1);
  assign w10[34] = |(datain[175:172] ^ 11);
  assign w10[35] = |(datain[171:168] ^ 4);
  assign w10[36] = |(datain[167:164] ^ 4);
  assign w10[37] = |(datain[163:160] ^ 0);
  assign w10[38] = |(datain[159:156] ^ 11);
  assign w10[39] = |(datain[155:152] ^ 9);
  assign w10[40] = |(datain[151:148] ^ 1);
  assign w10[41] = |(datain[147:144] ^ 6);
  assign w10[42] = |(datain[143:140] ^ 0);
  assign w10[43] = |(datain[139:136] ^ 9);
  assign w10[44] = |(datain[135:132] ^ 5);
  assign w10[45] = |(datain[131:128] ^ 10);
  assign w10[46] = |(datain[127:124] ^ 12);
  assign w10[47] = |(datain[123:120] ^ 13);
  assign w10[48] = |(datain[119:116] ^ 2);
  assign w10[49] = |(datain[115:112] ^ 1);
  assign w10[50] = |(datain[111:108] ^ 5);
  assign w10[51] = |(datain[107:104] ^ 15);
  assign w10[52] = |(datain[103:100] ^ 0);
  assign w10[53] = |(datain[99:96] ^ 7);
  assign w10[54] = |(datain[95:92] ^ 2);
  assign w10[55] = |(datain[91:88] ^ 6);
  assign w10[56] = |(datain[87:84] ^ 8);
  assign w10[57] = |(datain[83:80] ^ 0);
  assign w10[58] = |(datain[79:76] ^ 4);
  assign w10[59] = |(datain[75:72] ^ 13);
  assign w10[60] = |(datain[71:68] ^ 0);
  assign w10[61] = |(datain[67:64] ^ 6);
  assign w10[62] = |(datain[63:60] ^ 4);
  assign w10[63] = |(datain[59:56] ^ 0);
  assign w10[64] = |(datain[55:52] ^ 11);
  assign w10[65] = |(datain[51:48] ^ 4);
  assign w10[66] = |(datain[47:44] ^ 3);
  assign w10[67] = |(datain[43:40] ^ 14);
  assign w10[68] = |(datain[39:36] ^ 12);
  assign w10[69] = |(datain[35:32] ^ 13);
  assign w10[70] = |(datain[31:28] ^ 2);
  assign w10[71] = |(datain[27:24] ^ 1);
  assign w10[72] = |(datain[23:20] ^ 12);
  assign w10[73] = |(datain[19:16] ^ 3);
  assign comp[10] = ~(|w10);
  wire [76-1:0] w11;
  assign w11[0] = |(datain[311:308] ^ 0);
  assign w11[1] = |(datain[307:304] ^ 6);
  assign w11[2] = |(datain[303:300] ^ 8);
  assign w11[3] = |(datain[299:296] ^ 13);
  assign w11[4] = |(datain[295:292] ^ 11);
  assign w11[5] = |(datain[291:288] ^ 6);
  assign w11[6] = |(datain[287:284] ^ 0);
  assign w11[7] = |(datain[283:280] ^ 8);
  assign w11[8] = |(datain[279:276] ^ 0);
  assign w11[9] = |(datain[275:272] ^ 1);
  assign w11[10] = |(datain[271:268] ^ 14);
  assign w11[11] = |(datain[267:264] ^ 8);
  assign w11[12] = |(datain[263:260] ^ 6);
  assign w11[13] = |(datain[259:256] ^ 11);
  assign w11[14] = |(datain[255:252] ^ 0);
  assign w11[15] = |(datain[251:248] ^ 0);
  assign w11[16] = |(datain[247:244] ^ 5);
  assign w11[17] = |(datain[243:240] ^ 13);
  assign w11[18] = |(datain[239:236] ^ 5);
  assign w11[19] = |(datain[235:232] ^ 11);
  assign w11[20] = |(datain[231:228] ^ 8);
  assign w11[21] = |(datain[227:224] ^ 13);
  assign w11[22] = |(datain[223:220] ^ 9);
  assign w11[23] = |(datain[219:216] ^ 6);
  assign w11[24] = |(datain[215:212] ^ 10);
  assign w11[25] = |(datain[211:208] ^ 1);
  assign w11[26] = |(datain[207:204] ^ 0);
  assign w11[27] = |(datain[203:200] ^ 6);
  assign w11[28] = |(datain[199:196] ^ 11);
  assign w11[29] = |(datain[195:192] ^ 4);
  assign w11[30] = |(datain[191:188] ^ 4);
  assign w11[31] = |(datain[187:184] ^ 0);
  assign w11[32] = |(datain[183:180] ^ 12);
  assign w11[33] = |(datain[179:176] ^ 13);
  assign w11[34] = |(datain[175:172] ^ 2);
  assign w11[35] = |(datain[171:168] ^ 1);
  assign w11[36] = |(datain[167:164] ^ 8);
  assign w11[37] = |(datain[163:160] ^ 15);
  assign w11[38] = |(datain[159:156] ^ 8);
  assign w11[39] = |(datain[155:152] ^ 6);
  assign w11[40] = |(datain[151:148] ^ 0);
  assign w11[41] = |(datain[147:144] ^ 4);
  assign w11[42] = |(datain[143:140] ^ 0);
  assign w11[43] = |(datain[139:136] ^ 2);
  assign w11[44] = |(datain[135:132] ^ 11);
  assign w11[45] = |(datain[131:128] ^ 8);
  assign w11[46] = |(datain[127:124] ^ 0);
  assign w11[47] = |(datain[123:120] ^ 0);
  assign w11[48] = |(datain[119:116] ^ 4);
  assign w11[49] = |(datain[115:112] ^ 2);
  assign w11[50] = |(datain[111:108] ^ 14);
  assign w11[51] = |(datain[107:104] ^ 8);
  assign w11[52] = |(datain[103:100] ^ 2);
  assign w11[53] = |(datain[99:96] ^ 11);
  assign w11[54] = |(datain[95:92] ^ 0);
  assign w11[55] = |(datain[91:88] ^ 0);
  assign w11[56] = |(datain[87:84] ^ 8);
  assign w11[57] = |(datain[83:80] ^ 13);
  assign w11[58] = |(datain[79:76] ^ 9);
  assign w11[59] = |(datain[75:72] ^ 6);
  assign w11[60] = |(datain[71:68] ^ 15);
  assign w11[61] = |(datain[67:64] ^ 15);
  assign w11[62] = |(datain[63:60] ^ 0);
  assign w11[63] = |(datain[59:56] ^ 1);
  assign w11[64] = |(datain[55:52] ^ 11);
  assign w11[65] = |(datain[51:48] ^ 9);
  assign w11[66] = |(datain[47:44] ^ 0);
  assign w11[67] = |(datain[43:40] ^ 5);
  assign w11[68] = |(datain[39:36] ^ 0);
  assign w11[69] = |(datain[35:32] ^ 0);
  assign w11[70] = |(datain[31:28] ^ 11);
  assign w11[71] = |(datain[27:24] ^ 4);
  assign w11[72] = |(datain[23:20] ^ 4);
  assign w11[73] = |(datain[19:16] ^ 0);
  assign w11[74] = |(datain[15:12] ^ 12);
  assign w11[75] = |(datain[11:8] ^ 13);
  assign comp[11] = ~(|w11);
  wire [76-1:0] w12;
  assign w12[0] = |(datain[311:308] ^ 0);
  assign w12[1] = |(datain[307:304] ^ 4);
  assign w12[2] = |(datain[303:300] ^ 0);
  assign w12[3] = |(datain[299:296] ^ 2);
  assign w12[4] = |(datain[295:292] ^ 0);
  assign w12[5] = |(datain[291:288] ^ 5);
  assign w12[6] = |(datain[287:284] ^ 0);
  assign w12[7] = |(datain[283:280] ^ 2);
  assign w12[8] = |(datain[279:276] ^ 0);
  assign w12[9] = |(datain[275:272] ^ 0);
  assign w12[10] = |(datain[271:268] ^ 8);
  assign w12[11] = |(datain[267:264] ^ 9);
  assign w12[12] = |(datain[263:260] ^ 0);
  assign w12[13] = |(datain[259:256] ^ 4);
  assign w12[14] = |(datain[255:252] ^ 8);
  assign w12[15] = |(datain[251:248] ^ 13);
  assign w12[16] = |(datain[247:244] ^ 9);
  assign w12[17] = |(datain[243:240] ^ 6);
  assign w12[18] = |(datain[239:236] ^ 15);
  assign w12[19] = |(datain[235:232] ^ 10);
  assign w12[20] = |(datain[231:228] ^ 0);
  assign w12[21] = |(datain[227:224] ^ 1);
  assign w12[22] = |(datain[223:220] ^ 11);
  assign w12[23] = |(datain[219:216] ^ 9);
  assign w12[24] = |(datain[215:212] ^ 0);
  assign w12[25] = |(datain[211:208] ^ 5);
  assign w12[26] = |(datain[207:204] ^ 0);
  assign w12[27] = |(datain[203:200] ^ 0);
  assign w12[28] = |(datain[199:196] ^ 11);
  assign w12[29] = |(datain[195:192] ^ 4);
  assign w12[30] = |(datain[191:188] ^ 4);
  assign w12[31] = |(datain[187:184] ^ 0);
  assign w12[32] = |(datain[183:180] ^ 12);
  assign w12[33] = |(datain[179:176] ^ 13);
  assign w12[34] = |(datain[175:172] ^ 2);
  assign w12[35] = |(datain[171:168] ^ 1);
  assign w12[36] = |(datain[167:164] ^ 5);
  assign w12[37] = |(datain[163:160] ^ 3);
  assign w12[38] = |(datain[159:156] ^ 5);
  assign w12[39] = |(datain[155:152] ^ 5);
  assign w12[40] = |(datain[151:148] ^ 8);
  assign w12[41] = |(datain[147:144] ^ 11);
  assign w12[42] = |(datain[143:140] ^ 1);
  assign w12[43] = |(datain[139:136] ^ 4);
  assign w12[44] = |(datain[135:132] ^ 8);
  assign w12[45] = |(datain[131:128] ^ 1);
  assign w12[46] = |(datain[127:124] ^ 12);
  assign w12[47] = |(datain[123:120] ^ 2);
  assign w12[48] = |(datain[119:116] ^ 0);
  assign w12[49] = |(datain[115:112] ^ 3);
  assign w12[50] = |(datain[111:108] ^ 0);
  assign w12[51] = |(datain[107:104] ^ 1);
  assign w12[52] = |(datain[103:100] ^ 11);
  assign w12[53] = |(datain[99:96] ^ 9);
  assign w12[54] = |(datain[95:92] ^ 1);
  assign w12[55] = |(datain[91:88] ^ 9);
  assign w12[56] = |(datain[87:84] ^ 0);
  assign w12[57] = |(datain[83:80] ^ 5);
  assign w12[58] = |(datain[79:76] ^ 9);
  assign w12[59] = |(datain[75:72] ^ 0);
  assign w12[60] = |(datain[71:68] ^ 8);
  assign w12[61] = |(datain[67:64] ^ 13);
  assign w12[62] = |(datain[63:60] ^ 11);
  assign w12[63] = |(datain[59:56] ^ 14);
  assign w12[64] = |(datain[55:52] ^ 10);
  assign w12[65] = |(datain[51:48] ^ 1);
  assign w12[66] = |(datain[47:44] ^ 0);
  assign w12[67] = |(datain[43:40] ^ 6);
  assign w12[68] = |(datain[39:36] ^ 8);
  assign w12[69] = |(datain[35:32] ^ 13);
  assign w12[70] = |(datain[31:28] ^ 11);
  assign w12[71] = |(datain[27:24] ^ 6);
  assign w12[72] = |(datain[23:20] ^ 0);
  assign w12[73] = |(datain[19:16] ^ 8);
  assign w12[74] = |(datain[15:12] ^ 0);
  assign w12[75] = |(datain[11:8] ^ 1);
  assign comp[12] = ~(|w12);
  wire [74-1:0] w13;
  assign w13[0] = |(datain[311:308] ^ 8);
  assign w13[1] = |(datain[307:304] ^ 11);
  assign w13[2] = |(datain[303:300] ^ 13);
  assign w13[3] = |(datain[299:296] ^ 1);
  assign w13[4] = |(datain[295:292] ^ 11);
  assign w13[5] = |(datain[291:288] ^ 8);
  assign w13[6] = |(datain[287:284] ^ 0);
  assign w13[7] = |(datain[283:280] ^ 0);
  assign w13[8] = |(datain[279:276] ^ 4);
  assign w13[9] = |(datain[275:272] ^ 2);
  assign w13[10] = |(datain[271:268] ^ 12);
  assign w13[11] = |(datain[267:264] ^ 13);
  assign w13[12] = |(datain[263:260] ^ 2);
  assign w13[13] = |(datain[259:256] ^ 1);
  assign w13[14] = |(datain[255:252] ^ 5);
  assign w13[15] = |(datain[251:248] ^ 9);
  assign w13[16] = |(datain[247:244] ^ 0);
  assign w13[17] = |(datain[243:240] ^ 3);
  assign w13[18] = |(datain[239:236] ^ 0);
  assign w13[19] = |(datain[235:232] ^ 13);
  assign w13[20] = |(datain[231:228] ^ 11);
  assign w13[21] = |(datain[227:224] ^ 10);
  assign w13[22] = |(datain[223:220] ^ 0);
  assign w13[23] = |(datain[219:216] ^ 0);
  assign w13[24] = |(datain[215:212] ^ 0);
  assign w13[25] = |(datain[211:208] ^ 1);
  assign w13[26] = |(datain[207:204] ^ 11);
  assign w13[27] = |(datain[203:200] ^ 4);
  assign w13[28] = |(datain[199:196] ^ 4);
  assign w13[29] = |(datain[195:192] ^ 0);
  assign w13[30] = |(datain[191:188] ^ 12);
  assign w13[31] = |(datain[187:184] ^ 13);
  assign w13[32] = |(datain[183:180] ^ 2);
  assign w13[33] = |(datain[179:176] ^ 1);
  assign w13[34] = |(datain[175:172] ^ 1);
  assign w13[35] = |(datain[171:168] ^ 15);
  assign w13[36] = |(datain[167:164] ^ 11);
  assign w13[37] = |(datain[163:160] ^ 8);
  assign w13[38] = |(datain[159:156] ^ 0);
  assign w13[39] = |(datain[155:152] ^ 0);
  assign w13[40] = |(datain[151:148] ^ 5);
  assign w13[41] = |(datain[147:144] ^ 7);
  assign w13[42] = |(datain[143:140] ^ 12);
  assign w13[43] = |(datain[139:136] ^ 13);
  assign w13[44] = |(datain[135:132] ^ 2);
  assign w13[45] = |(datain[131:128] ^ 1);
  assign w13[46] = |(datain[127:124] ^ 5);
  assign w13[47] = |(datain[123:120] ^ 2);
  assign w13[48] = |(datain[119:116] ^ 8);
  assign w13[49] = |(datain[115:112] ^ 11);
  assign w13[50] = |(datain[111:108] ^ 12);
  assign w13[51] = |(datain[107:104] ^ 1);
  assign w13[52] = |(datain[103:100] ^ 3);
  assign w13[53] = |(datain[99:96] ^ 3);
  assign w13[54] = |(datain[95:92] ^ 12);
  assign w13[55] = |(datain[91:88] ^ 2);
  assign w13[56] = |(datain[87:84] ^ 11);
  assign w13[57] = |(datain[83:80] ^ 9);
  assign w13[58] = |(datain[79:76] ^ 0);
  assign w13[59] = |(datain[75:72] ^ 10);
  assign w13[60] = |(datain[71:68] ^ 0);
  assign w13[61] = |(datain[67:64] ^ 0);
  assign w13[62] = |(datain[63:60] ^ 3);
  assign w13[63] = |(datain[59:56] ^ 3);
  assign w13[64] = |(datain[55:52] ^ 13);
  assign w13[65] = |(datain[51:48] ^ 2);
  assign w13[66] = |(datain[47:44] ^ 15);
  assign w13[67] = |(datain[43:40] ^ 7);
  assign w13[68] = |(datain[39:36] ^ 15);
  assign w13[69] = |(datain[35:32] ^ 1);
  assign w13[70] = |(datain[31:28] ^ 15);
  assign w13[71] = |(datain[27:24] ^ 7);
  assign w13[72] = |(datain[23:20] ^ 14);
  assign w13[73] = |(datain[19:16] ^ 1);
  assign comp[13] = ~(|w13);
  wire [74-1:0] w14;
  assign w14[0] = |(datain[311:308] ^ 14);
  assign w14[1] = |(datain[307:304] ^ 8);
  assign w14[2] = |(datain[303:300] ^ 10);
  assign w14[3] = |(datain[299:296] ^ 15);
  assign w14[4] = |(datain[295:292] ^ 0);
  assign w14[5] = |(datain[291:288] ^ 0);
  assign w14[6] = |(datain[287:284] ^ 5);
  assign w14[7] = |(datain[283:280] ^ 11);
  assign w14[8] = |(datain[279:276] ^ 5);
  assign w14[9] = |(datain[275:272] ^ 8);
  assign w14[10] = |(datain[271:268] ^ 0);
  assign w14[11] = |(datain[267:264] ^ 3);
  assign w14[12] = |(datain[263:260] ^ 12);
  assign w14[13] = |(datain[259:256] ^ 1);
  assign w14[14] = |(datain[255:252] ^ 15);
  assign w14[15] = |(datain[251:248] ^ 7);
  assign w14[16] = |(datain[247:244] ^ 13);
  assign w14[17] = |(datain[243:240] ^ 8);
  assign w14[18] = |(datain[239:236] ^ 3);
  assign w14[19] = |(datain[235:232] ^ 2);
  assign w14[20] = |(datain[231:228] ^ 14);
  assign w14[21] = |(datain[227:224] ^ 4);
  assign w14[22] = |(datain[223:220] ^ 0);
  assign w14[23] = |(datain[219:216] ^ 3);
  assign w14[24] = |(datain[215:212] ^ 12);
  assign w14[25] = |(datain[211:208] ^ 8);
  assign w14[26] = |(datain[207:204] ^ 11);
  assign w14[27] = |(datain[203:200] ^ 4);
  assign w14[28] = |(datain[199:196] ^ 4);
  assign w14[29] = |(datain[195:192] ^ 0);
  assign w14[30] = |(datain[191:188] ^ 12);
  assign w14[31] = |(datain[187:184] ^ 13);
  assign w14[32] = |(datain[183:180] ^ 2);
  assign w14[33] = |(datain[179:176] ^ 1);
  assign w14[34] = |(datain[175:172] ^ 0);
  assign w14[35] = |(datain[171:168] ^ 14);
  assign w14[36] = |(datain[167:164] ^ 1);
  assign w14[37] = |(datain[163:160] ^ 15);
  assign w14[38] = |(datain[159:156] ^ 7);
  assign w14[39] = |(datain[155:152] ^ 2);
  assign w14[40] = |(datain[151:148] ^ 1);
  assign w14[41] = |(datain[147:144] ^ 5);
  assign w14[42] = |(datain[143:140] ^ 2);
  assign w14[43] = |(datain[139:136] ^ 11);
  assign w14[44] = |(datain[135:132] ^ 12);
  assign w14[45] = |(datain[131:128] ^ 8);
  assign w14[46] = |(datain[127:124] ^ 7);
  assign w14[47] = |(datain[123:120] ^ 5);
  assign w14[48] = |(datain[119:116] ^ 1);
  assign w14[49] = |(datain[115:112] ^ 1);
  assign w14[50] = |(datain[111:108] ^ 3);
  assign w14[51] = |(datain[107:104] ^ 3);
  assign w14[52] = |(datain[103:100] ^ 13);
  assign w14[53] = |(datain[99:96] ^ 2);
  assign w14[54] = |(datain[95:92] ^ 11);
  assign w14[55] = |(datain[91:88] ^ 8);
  assign w14[56] = |(datain[87:84] ^ 0);
  assign w14[57] = |(datain[83:80] ^ 0);
  assign w14[58] = |(datain[79:76] ^ 4);
  assign w14[59] = |(datain[75:72] ^ 2);
  assign w14[60] = |(datain[71:68] ^ 12);
  assign w14[61] = |(datain[67:64] ^ 13);
  assign w14[62] = |(datain[63:60] ^ 2);
  assign w14[63] = |(datain[59:56] ^ 1);
  assign w14[64] = |(datain[55:52] ^ 11);
  assign w14[65] = |(datain[51:48] ^ 10);
  assign w14[66] = |(datain[47:44] ^ 9);
  assign w14[67] = |(datain[43:40] ^ 11);
  assign w14[68] = |(datain[39:36] ^ 0);
  assign w14[69] = |(datain[35:32] ^ 2);
  assign w14[70] = |(datain[31:28] ^ 11);
  assign w14[71] = |(datain[27:24] ^ 9);
  assign w14[72] = |(datain[23:20] ^ 0);
  assign w14[73] = |(datain[19:16] ^ 3);
  assign comp[14] = ~(|w14);
  wire [74-1:0] w15;
  assign w15[0] = |(datain[311:308] ^ 3);
  assign w15[1] = |(datain[307:304] ^ 3);
  assign w15[2] = |(datain[303:300] ^ 13);
  assign w15[3] = |(datain[299:296] ^ 2);
  assign w15[4] = |(datain[295:292] ^ 11);
  assign w15[5] = |(datain[291:288] ^ 8);
  assign w15[6] = |(datain[287:284] ^ 0);
  assign w15[7] = |(datain[283:280] ^ 0);
  assign w15[8] = |(datain[279:276] ^ 4);
  assign w15[9] = |(datain[275:272] ^ 2);
  assign w15[10] = |(datain[271:268] ^ 12);
  assign w15[11] = |(datain[267:264] ^ 13);
  assign w15[12] = |(datain[263:260] ^ 2);
  assign w15[13] = |(datain[259:256] ^ 1);
  assign w15[14] = |(datain[255:252] ^ 11);
  assign w15[15] = |(datain[251:248] ^ 10);
  assign w15[16] = |(datain[247:244] ^ 9);
  assign w15[17] = |(datain[243:240] ^ 11);
  assign w15[18] = |(datain[239:236] ^ 0);
  assign w15[19] = |(datain[235:232] ^ 2);
  assign w15[20] = |(datain[231:228] ^ 11);
  assign w15[21] = |(datain[227:224] ^ 9);
  assign w15[22] = |(datain[223:220] ^ 0);
  assign w15[23] = |(datain[219:216] ^ 3);
  assign w15[24] = |(datain[215:212] ^ 0);
  assign w15[25] = |(datain[211:208] ^ 0);
  assign w15[26] = |(datain[207:204] ^ 11);
  assign w15[27] = |(datain[203:200] ^ 4);
  assign w15[28] = |(datain[199:196] ^ 4);
  assign w15[29] = |(datain[195:192] ^ 0);
  assign w15[30] = |(datain[191:188] ^ 12);
  assign w15[31] = |(datain[187:184] ^ 13);
  assign w15[32] = |(datain[183:180] ^ 2);
  assign w15[33] = |(datain[179:176] ^ 1);
  assign w15[34] = |(datain[175:172] ^ 5);
  assign w15[35] = |(datain[171:168] ^ 9);
  assign w15[36] = |(datain[167:164] ^ 5);
  assign w15[37] = |(datain[163:160] ^ 10);
  assign w15[38] = |(datain[159:156] ^ 11);
  assign w15[39] = |(datain[155:152] ^ 8);
  assign w15[40] = |(datain[151:148] ^ 0);
  assign w15[41] = |(datain[147:144] ^ 1);
  assign w15[42] = |(datain[143:140] ^ 5);
  assign w15[43] = |(datain[139:136] ^ 7);
  assign w15[44] = |(datain[135:132] ^ 12);
  assign w15[45] = |(datain[131:128] ^ 13);
  assign w15[46] = |(datain[127:124] ^ 2);
  assign w15[47] = |(datain[123:120] ^ 1);
  assign w15[48] = |(datain[119:116] ^ 11);
  assign w15[49] = |(datain[115:112] ^ 4);
  assign w15[50] = |(datain[111:108] ^ 3);
  assign w15[51] = |(datain[107:104] ^ 14);
  assign w15[52] = |(datain[103:100] ^ 12);
  assign w15[53] = |(datain[99:96] ^ 13);
  assign w15[54] = |(datain[95:92] ^ 2);
  assign w15[55] = |(datain[91:88] ^ 1);
  assign w15[56] = |(datain[87:84] ^ 14);
  assign w15[57] = |(datain[83:80] ^ 9);
  assign w15[58] = |(datain[79:76] ^ 2);
  assign w15[59] = |(datain[75:72] ^ 12);
  assign w15[60] = |(datain[71:68] ^ 15);
  assign w15[61] = |(datain[67:64] ^ 15);
  assign w15[62] = |(datain[63:60] ^ 11);
  assign w15[63] = |(datain[59:56] ^ 0);
  assign w15[64] = |(datain[55:52] ^ 0);
  assign w15[65] = |(datain[51:48] ^ 3);
  assign w15[66] = |(datain[47:44] ^ 12);
  assign w15[67] = |(datain[43:40] ^ 15);
  assign w15[68] = |(datain[39:36] ^ 2);
  assign w15[69] = |(datain[35:32] ^ 10);
  assign w15[70] = |(datain[31:28] ^ 2);
  assign w15[71] = |(datain[27:24] ^ 14);
  assign w15[72] = |(datain[23:20] ^ 2);
  assign w15[73] = |(datain[19:16] ^ 10);
  assign comp[15] = ~(|w15);
  wire [74-1:0] w16;
  assign w16[0] = |(datain[311:308] ^ 5);
  assign w16[1] = |(datain[307:304] ^ 8);
  assign w16[2] = |(datain[303:300] ^ 8);
  assign w16[3] = |(datain[299:296] ^ 0);
  assign w16[4] = |(datain[295:292] ^ 15);
  assign w16[5] = |(datain[291:288] ^ 12);
  assign w16[6] = |(datain[287:284] ^ 0);
  assign w16[7] = |(datain[283:280] ^ 0);
  assign w16[8] = |(datain[279:276] ^ 7);
  assign w16[9] = |(datain[275:272] ^ 4);
  assign w16[10] = |(datain[271:268] ^ 1);
  assign w16[11] = |(datain[267:264] ^ 4);
  assign w16[12] = |(datain[263:260] ^ 8);
  assign w16[13] = |(datain[259:256] ^ 10);
  assign w16[14] = |(datain[255:252] ^ 12);
  assign w16[15] = |(datain[251:248] ^ 12);
  assign w16[16] = |(datain[247:244] ^ 3);
  assign w16[17] = |(datain[243:240] ^ 2);
  assign w16[18] = |(datain[239:236] ^ 14);
  assign w16[19] = |(datain[235:232] ^ 13);
  assign w16[20] = |(datain[231:228] ^ 11);
  assign w16[21] = |(datain[227:224] ^ 4);
  assign w16[22] = |(datain[223:220] ^ 4);
  assign w16[23] = |(datain[219:216] ^ 0);
  assign w16[24] = |(datain[215:212] ^ 1);
  assign w16[25] = |(datain[211:208] ^ 14);
  assign w16[26] = |(datain[207:204] ^ 0);
  assign w16[27] = |(datain[203:200] ^ 6);
  assign w16[28] = |(datain[199:196] ^ 1);
  assign w16[29] = |(datain[195:192] ^ 15);
  assign w16[30] = |(datain[191:188] ^ 12);
  assign w16[31] = |(datain[187:184] ^ 13);
  assign w16[32] = |(datain[183:180] ^ 2);
  assign w16[33] = |(datain[179:176] ^ 1);
  assign w16[34] = |(datain[175:172] ^ 1);
  assign w16[35] = |(datain[171:168] ^ 15);
  assign w16[36] = |(datain[167:164] ^ 7);
  assign w16[37] = |(datain[163:160] ^ 3);
  assign w16[38] = |(datain[159:156] ^ 0);
  assign w16[39] = |(datain[155:152] ^ 6);
  assign w16[40] = |(datain[151:148] ^ 14);
  assign w16[41] = |(datain[147:144] ^ 8);
  assign w16[42] = |(datain[143:140] ^ 6);
  assign w16[43] = |(datain[139:136] ^ 14);
  assign w16[44] = |(datain[135:132] ^ 0);
  assign w16[45] = |(datain[131:128] ^ 0);
  assign w16[46] = |(datain[127:124] ^ 14);
  assign w16[47] = |(datain[123:120] ^ 11);
  assign w16[48] = |(datain[119:116] ^ 2);
  assign w16[49] = |(datain[115:112] ^ 4);
  assign w16[50] = |(datain[111:108] ^ 9);
  assign w16[51] = |(datain[107:104] ^ 0);
  assign w16[52] = |(datain[103:100] ^ 0);
  assign w16[53] = |(datain[99:96] ^ 14);
  assign w16[54] = |(datain[95:92] ^ 1);
  assign w16[55] = |(datain[91:88] ^ 15);
  assign w16[56] = |(datain[87:84] ^ 11);
  assign w16[57] = |(datain[83:80] ^ 8);
  assign w16[58] = |(datain[79:76] ^ 0);
  assign w16[59] = |(datain[75:72] ^ 0);
  assign w16[60] = |(datain[71:68] ^ 4);
  assign w16[61] = |(datain[67:64] ^ 2);
  assign w16[62] = |(datain[63:60] ^ 3);
  assign w16[63] = |(datain[59:56] ^ 3);
  assign w16[64] = |(datain[55:52] ^ 12);
  assign w16[65] = |(datain[51:48] ^ 9);
  assign w16[66] = |(datain[47:44] ^ 3);
  assign w16[67] = |(datain[43:40] ^ 3);
  assign w16[68] = |(datain[39:36] ^ 13);
  assign w16[69] = |(datain[35:32] ^ 2);
  assign w16[70] = |(datain[31:28] ^ 12);
  assign w16[71] = |(datain[27:24] ^ 13);
  assign w16[72] = |(datain[23:20] ^ 2);
  assign w16[73] = |(datain[19:16] ^ 1);
  assign comp[16] = ~(|w16);
  wire [74-1:0] w17;
  assign w17[0] = |(datain[311:308] ^ 3);
  assign w17[1] = |(datain[307:304] ^ 3);
  assign w17[2] = |(datain[303:300] ^ 12);
  assign w17[3] = |(datain[299:296] ^ 9);
  assign w17[4] = |(datain[295:292] ^ 3);
  assign w17[5] = |(datain[291:288] ^ 3);
  assign w17[6] = |(datain[287:284] ^ 13);
  assign w17[7] = |(datain[283:280] ^ 2);
  assign w17[8] = |(datain[279:276] ^ 12);
  assign w17[9] = |(datain[275:272] ^ 13);
  assign w17[10] = |(datain[271:268] ^ 2);
  assign w17[11] = |(datain[267:264] ^ 1);
  assign w17[12] = |(datain[263:260] ^ 11);
  assign w17[13] = |(datain[259:256] ^ 4);
  assign w17[14] = |(datain[255:252] ^ 4);
  assign w17[15] = |(datain[251:248] ^ 0);
  assign w17[16] = |(datain[247:244] ^ 8);
  assign w17[17] = |(datain[243:240] ^ 13);
  assign w17[18] = |(datain[239:236] ^ 9);
  assign w17[19] = |(datain[235:232] ^ 6);
  assign w17[20] = |(datain[231:228] ^ 7);
  assign w17[21] = |(datain[227:224] ^ 6);
  assign w17[22] = |(datain[223:220] ^ 0);
  assign w17[23] = |(datain[219:216] ^ 4);
  assign w17[24] = |(datain[215:212] ^ 11);
  assign w17[25] = |(datain[211:208] ^ 9);
  assign w17[26] = |(datain[207:204] ^ 0);
  assign w17[27] = |(datain[203:200] ^ 3);
  assign w17[28] = |(datain[199:196] ^ 0);
  assign w17[29] = |(datain[195:192] ^ 0);
  assign w17[30] = |(datain[191:188] ^ 12);
  assign w17[31] = |(datain[187:184] ^ 13);
  assign w17[32] = |(datain[183:180] ^ 2);
  assign w17[33] = |(datain[179:176] ^ 1);
  assign w17[34] = |(datain[175:172] ^ 10);
  assign w17[35] = |(datain[171:168] ^ 1);
  assign w17[36] = |(datain[167:164] ^ 9);
  assign w17[37] = |(datain[163:160] ^ 6);
  assign w17[38] = |(datain[159:156] ^ 0);
  assign w17[39] = |(datain[155:152] ^ 0);
  assign w17[40] = |(datain[151:148] ^ 2);
  assign w17[41] = |(datain[147:144] ^ 4);
  assign w17[42] = |(datain[143:140] ^ 14);
  assign w17[43] = |(datain[139:136] ^ 0);
  assign w17[44] = |(datain[135:132] ^ 0);
  assign w17[45] = |(datain[131:128] ^ 12);
  assign w17[46] = |(datain[127:124] ^ 0);
  assign w17[47] = |(datain[123:120] ^ 12);
  assign w17[48] = |(datain[119:116] ^ 10);
  assign w17[49] = |(datain[115:112] ^ 3);
  assign w17[50] = |(datain[111:108] ^ 9);
  assign w17[51] = |(datain[107:104] ^ 6);
  assign w17[52] = |(datain[103:100] ^ 0);
  assign w17[53] = |(datain[99:96] ^ 0);
  assign w17[54] = |(datain[95:92] ^ 14);
  assign w17[55] = |(datain[91:88] ^ 8);
  assign w17[56] = |(datain[87:84] ^ 4);
  assign w17[57] = |(datain[83:80] ^ 8);
  assign w17[58] = |(datain[79:76] ^ 0);
  assign w17[59] = |(datain[75:72] ^ 0);
  assign w17[60] = |(datain[71:68] ^ 0);
  assign w17[61] = |(datain[67:64] ^ 6);
  assign w17[62] = |(datain[63:60] ^ 3);
  assign w17[63] = |(datain[59:56] ^ 3);
  assign w17[64] = |(datain[55:52] ^ 12);
  assign w17[65] = |(datain[51:48] ^ 0);
  assign w17[66] = |(datain[47:44] ^ 8);
  assign w17[67] = |(datain[43:40] ^ 14);
  assign w17[68] = |(datain[39:36] ^ 12);
  assign w17[69] = |(datain[35:32] ^ 0);
  assign w17[70] = |(datain[31:28] ^ 15);
  assign w17[71] = |(datain[27:24] ^ 10);
  assign w17[72] = |(datain[23:20] ^ 10);
  assign w17[73] = |(datain[19:16] ^ 1);
  assign comp[17] = ~(|w17);
  wire [74-1:0] w18;
  assign w18[0] = |(datain[311:308] ^ 3);
  assign w18[1] = |(datain[307:304] ^ 3);
  assign w18[2] = |(datain[303:300] ^ 15);
  assign w18[3] = |(datain[299:296] ^ 6);
  assign w18[4] = |(datain[295:292] ^ 8);
  assign w18[5] = |(datain[291:288] ^ 1);
  assign w18[6] = |(datain[287:284] ^ 12);
  assign w18[7] = |(datain[283:280] ^ 5);
  assign w18[8] = |(datain[279:276] ^ 0);
  assign w18[9] = |(datain[275:272] ^ 0);
  assign w18[10] = |(datain[271:268] ^ 0);
  assign w18[11] = |(datain[267:264] ^ 1);
  assign w18[12] = |(datain[263:260] ^ 14);
  assign w18[13] = |(datain[259:256] ^ 8);
  assign w18[14] = |(datain[255:252] ^ 8);
  assign w18[15] = |(datain[251:248] ^ 7);
  assign w18[16] = |(datain[247:244] ^ 0);
  assign w18[17] = |(datain[243:240] ^ 1);
  assign w18[18] = |(datain[239:236] ^ 11);
  assign w18[19] = |(datain[235:232] ^ 4);
  assign w18[20] = |(datain[231:228] ^ 4);
  assign w18[21] = |(datain[227:224] ^ 0);
  assign w18[22] = |(datain[223:220] ^ 11);
  assign w18[23] = |(datain[219:216] ^ 9);
  assign w18[24] = |(datain[215:212] ^ 12);
  assign w18[25] = |(datain[211:208] ^ 1);
  assign w18[26] = |(datain[207:204] ^ 0);
  assign w18[27] = |(datain[203:200] ^ 4);
  assign w18[28] = |(datain[199:196] ^ 5);
  assign w18[29] = |(datain[195:192] ^ 10);
  assign w18[30] = |(datain[191:188] ^ 12);
  assign w18[31] = |(datain[187:184] ^ 13);
  assign w18[32] = |(datain[183:180] ^ 2);
  assign w18[33] = |(datain[179:176] ^ 1);
  assign w18[34] = |(datain[175:172] ^ 11);
  assign w18[35] = |(datain[171:168] ^ 8);
  assign w18[36] = |(datain[167:164] ^ 0);
  assign w18[37] = |(datain[163:160] ^ 0);
  assign w18[38] = |(datain[159:156] ^ 4);
  assign w18[39] = |(datain[155:152] ^ 2);
  assign w18[40] = |(datain[151:148] ^ 14);
  assign w18[41] = |(datain[147:144] ^ 8);
  assign w18[42] = |(datain[143:140] ^ 4);
  assign w18[43] = |(datain[139:136] ^ 0);
  assign w18[44] = |(datain[135:132] ^ 0);
  assign w18[45] = |(datain[131:128] ^ 0);
  assign w18[46] = |(datain[127:124] ^ 11);
  assign w18[47] = |(datain[123:120] ^ 4);
  assign w18[48] = |(datain[119:116] ^ 4);
  assign w18[49] = |(datain[115:112] ^ 0);
  assign w18[50] = |(datain[111:108] ^ 11);
  assign w18[51] = |(datain[107:104] ^ 9);
  assign w18[52] = |(datain[103:100] ^ 0);
  assign w18[53] = |(datain[99:96] ^ 4);
  assign w18[54] = |(datain[95:92] ^ 0);
  assign w18[55] = |(datain[91:88] ^ 0);
  assign w18[56] = |(datain[87:84] ^ 11);
  assign w18[57] = |(datain[83:80] ^ 10);
  assign w18[58] = |(datain[79:76] ^ 2);
  assign w18[59] = |(datain[75:72] ^ 0);
  assign w18[60] = |(datain[71:68] ^ 0);
  assign w18[61] = |(datain[67:64] ^ 3);
  assign w18[62] = |(datain[63:60] ^ 12);
  assign w18[63] = |(datain[59:56] ^ 13);
  assign w18[64] = |(datain[55:52] ^ 2);
  assign w18[65] = |(datain[51:48] ^ 1);
  assign w18[66] = |(datain[47:44] ^ 11);
  assign w18[67] = |(datain[43:40] ^ 8);
  assign w18[68] = |(datain[39:36] ^ 0);
  assign w18[69] = |(datain[35:32] ^ 1);
  assign w18[70] = |(datain[31:28] ^ 5);
  assign w18[71] = |(datain[27:24] ^ 7);
  assign w18[72] = |(datain[23:20] ^ 2);
  assign w18[73] = |(datain[19:16] ^ 14);
  assign comp[18] = ~(|w18);
  wire [74-1:0] w19;
  assign w19[0] = |(datain[311:308] ^ 2);
  assign w19[1] = |(datain[307:304] ^ 1);
  assign w19[2] = |(datain[303:300] ^ 11);
  assign w19[3] = |(datain[299:296] ^ 8);
  assign w19[4] = |(datain[295:292] ^ 0);
  assign w19[5] = |(datain[291:288] ^ 0);
  assign w19[6] = |(datain[287:284] ^ 4);
  assign w19[7] = |(datain[283:280] ^ 2);
  assign w19[8] = |(datain[279:276] ^ 14);
  assign w19[9] = |(datain[275:272] ^ 8);
  assign w19[10] = |(datain[271:268] ^ 4);
  assign w19[11] = |(datain[267:264] ^ 0);
  assign w19[12] = |(datain[263:260] ^ 0);
  assign w19[13] = |(datain[259:256] ^ 0);
  assign w19[14] = |(datain[255:252] ^ 11);
  assign w19[15] = |(datain[251:248] ^ 4);
  assign w19[16] = |(datain[247:244] ^ 4);
  assign w19[17] = |(datain[243:240] ^ 0);
  assign w19[18] = |(datain[239:236] ^ 11);
  assign w19[19] = |(datain[235:232] ^ 9);
  assign w19[20] = |(datain[231:228] ^ 0);
  assign w19[21] = |(datain[227:224] ^ 4);
  assign w19[22] = |(datain[223:220] ^ 0);
  assign w19[23] = |(datain[219:216] ^ 0);
  assign w19[24] = |(datain[215:212] ^ 11);
  assign w19[25] = |(datain[211:208] ^ 10);
  assign w19[26] = |(datain[207:204] ^ 2);
  assign w19[27] = |(datain[203:200] ^ 0);
  assign w19[28] = |(datain[199:196] ^ 0);
  assign w19[29] = |(datain[195:192] ^ 3);
  assign w19[30] = |(datain[191:188] ^ 12);
  assign w19[31] = |(datain[187:184] ^ 13);
  assign w19[32] = |(datain[183:180] ^ 2);
  assign w19[33] = |(datain[179:176] ^ 1);
  assign w19[34] = |(datain[175:172] ^ 11);
  assign w19[35] = |(datain[171:168] ^ 8);
  assign w19[36] = |(datain[167:164] ^ 0);
  assign w19[37] = |(datain[163:160] ^ 1);
  assign w19[38] = |(datain[159:156] ^ 5);
  assign w19[39] = |(datain[155:152] ^ 7);
  assign w19[40] = |(datain[151:148] ^ 2);
  assign w19[41] = |(datain[147:144] ^ 14);
  assign w19[42] = |(datain[143:140] ^ 8);
  assign w19[43] = |(datain[139:136] ^ 11);
  assign w19[44] = |(datain[135:132] ^ 1);
  assign w19[45] = |(datain[131:128] ^ 6);
  assign w19[46] = |(datain[127:124] ^ 1);
  assign w19[47] = |(datain[123:120] ^ 2);
  assign w19[48] = |(datain[119:116] ^ 0);
  assign w19[49] = |(datain[115:112] ^ 3);
  assign w19[50] = |(datain[111:108] ^ 2);
  assign w19[51] = |(datain[107:104] ^ 14);
  assign w19[52] = |(datain[103:100] ^ 8);
  assign w19[53] = |(datain[99:96] ^ 11);
  assign w19[54] = |(datain[95:92] ^ 0);
  assign w19[55] = |(datain[91:88] ^ 14);
  assign w19[56] = |(datain[87:84] ^ 1);
  assign w19[57] = |(datain[83:80] ^ 0);
  assign w19[58] = |(datain[79:76] ^ 0);
  assign w19[59] = |(datain[75:72] ^ 3);
  assign w19[60] = |(datain[71:68] ^ 8);
  assign w19[61] = |(datain[67:64] ^ 0);
  assign w19[62] = |(datain[63:60] ^ 14);
  assign w19[63] = |(datain[59:56] ^ 1);
  assign w19[64] = |(datain[55:52] ^ 14);
  assign w19[65] = |(datain[51:48] ^ 0);
  assign w19[66] = |(datain[47:44] ^ 15);
  assign w19[67] = |(datain[43:40] ^ 14);
  assign w19[68] = |(datain[39:36] ^ 12);
  assign w19[69] = |(datain[35:32] ^ 1);
  assign w19[70] = |(datain[31:28] ^ 12);
  assign w19[71] = |(datain[27:24] ^ 13);
  assign w19[72] = |(datain[23:20] ^ 2);
  assign w19[73] = |(datain[19:16] ^ 1);
  assign comp[19] = ~(|w19);
  wire [74-1:0] w20;
  assign w20[0] = |(datain[311:308] ^ 11);
  assign w20[1] = |(datain[307:304] ^ 4);
  assign w20[2] = |(datain[303:300] ^ 4);
  assign w20[3] = |(datain[299:296] ^ 0);
  assign w20[4] = |(datain[295:292] ^ 8);
  assign w20[5] = |(datain[291:288] ^ 13);
  assign w20[6] = |(datain[287:284] ^ 9);
  assign w20[7] = |(datain[283:280] ^ 6);
  assign w20[8] = |(datain[279:276] ^ 14);
  assign w20[9] = |(datain[275:272] ^ 15);
  assign w20[10] = |(datain[271:268] ^ 0);
  assign w20[11] = |(datain[267:264] ^ 4);
  assign w20[12] = |(datain[263:260] ^ 12);
  assign w20[13] = |(datain[259:256] ^ 13);
  assign w20[14] = |(datain[255:252] ^ 2);
  assign w20[15] = |(datain[251:248] ^ 1);
  assign w20[16] = |(datain[247:244] ^ 11);
  assign w20[17] = |(datain[243:240] ^ 4);
  assign w20[18] = |(datain[239:236] ^ 4);
  assign w20[19] = |(datain[235:232] ^ 0);
  assign w20[20] = |(datain[231:228] ^ 5);
  assign w20[21] = |(datain[227:224] ^ 9);
  assign w20[22] = |(datain[223:220] ^ 8);
  assign w20[23] = |(datain[219:216] ^ 13);
  assign w20[24] = |(datain[215:212] ^ 9);
  assign w20[25] = |(datain[211:208] ^ 6);
  assign w20[26] = |(datain[207:204] ^ 8);
  assign w20[27] = |(datain[203:200] ^ 11);
  assign w20[28] = |(datain[199:196] ^ 0);
  assign w20[29] = |(datain[195:192] ^ 5);
  assign w20[30] = |(datain[191:188] ^ 12);
  assign w20[31] = |(datain[187:184] ^ 13);
  assign w20[32] = |(datain[183:180] ^ 2);
  assign w20[33] = |(datain[179:176] ^ 1);
  assign w20[34] = |(datain[175:172] ^ 3);
  assign w20[35] = |(datain[171:168] ^ 2);
  assign w20[36] = |(datain[167:164] ^ 12);
  assign w20[37] = |(datain[163:160] ^ 0);
  assign w20[38] = |(datain[159:156] ^ 14);
  assign w20[39] = |(datain[155:152] ^ 8);
  assign w20[40] = |(datain[151:148] ^ 2);
  assign w20[41] = |(datain[147:144] ^ 9);
  assign w20[42] = |(datain[143:140] ^ 0);
  assign w20[43] = |(datain[139:136] ^ 0);
  assign w20[44] = |(datain[135:132] ^ 8);
  assign w20[45] = |(datain[131:128] ^ 13);
  assign w20[46] = |(datain[127:124] ^ 9);
  assign w20[47] = |(datain[123:120] ^ 6);
  assign w20[48] = |(datain[119:116] ^ 14);
  assign w20[49] = |(datain[115:112] ^ 11);
  assign w20[50] = |(datain[111:108] ^ 0);
  assign w20[51] = |(datain[107:104] ^ 4);
  assign w20[52] = |(datain[103:100] ^ 12);
  assign w20[53] = |(datain[99:96] ^ 13);
  assign w20[54] = |(datain[95:92] ^ 2);
  assign w20[55] = |(datain[91:88] ^ 1);
  assign w20[56] = |(datain[87:84] ^ 5);
  assign w20[57] = |(datain[83:80] ^ 10);
  assign w20[58] = |(datain[79:76] ^ 5);
  assign w20[59] = |(datain[75:72] ^ 9);
  assign w20[60] = |(datain[71:68] ^ 8);
  assign w20[61] = |(datain[67:64] ^ 0);
  assign w20[62] = |(datain[63:60] ^ 14);
  assign w20[63] = |(datain[59:56] ^ 1);
  assign w20[64] = |(datain[55:52] ^ 14);
  assign w20[65] = |(datain[51:48] ^ 0);
  assign w20[66] = |(datain[47:44] ^ 8);
  assign w20[67] = |(datain[43:40] ^ 0);
  assign w20[68] = |(datain[39:36] ^ 12);
  assign w20[69] = |(datain[35:32] ^ 9);
  assign w20[70] = |(datain[31:28] ^ 1);
  assign w20[71] = |(datain[27:24] ^ 15);
  assign w20[72] = |(datain[23:20] ^ 11);
  assign w20[73] = |(datain[19:16] ^ 8);
  assign comp[20] = ~(|w20);
  wire [76-1:0] w21;
  assign w21[0] = |(datain[311:308] ^ 5);
  assign w21[1] = |(datain[307:304] ^ 9);
  assign w21[2] = |(datain[303:300] ^ 8);
  assign w21[3] = |(datain[299:296] ^ 13);
  assign w21[4] = |(datain[295:292] ^ 9);
  assign w21[5] = |(datain[291:288] ^ 6);
  assign w21[6] = |(datain[287:284] ^ 8);
  assign w21[7] = |(datain[283:280] ^ 11);
  assign w21[8] = |(datain[279:276] ^ 0);
  assign w21[9] = |(datain[275:272] ^ 5);
  assign w21[10] = |(datain[271:268] ^ 12);
  assign w21[11] = |(datain[267:264] ^ 13);
  assign w21[12] = |(datain[263:260] ^ 2);
  assign w21[13] = |(datain[259:256] ^ 1);
  assign w21[14] = |(datain[255:252] ^ 3);
  assign w21[15] = |(datain[251:248] ^ 2);
  assign w21[16] = |(datain[247:244] ^ 12);
  assign w21[17] = |(datain[243:240] ^ 0);
  assign w21[18] = |(datain[239:236] ^ 14);
  assign w21[19] = |(datain[235:232] ^ 8);
  assign w21[20] = |(datain[231:228] ^ 2);
  assign w21[21] = |(datain[227:224] ^ 9);
  assign w21[22] = |(datain[223:220] ^ 0);
  assign w21[23] = |(datain[219:216] ^ 0);
  assign w21[24] = |(datain[215:212] ^ 8);
  assign w21[25] = |(datain[211:208] ^ 13);
  assign w21[26] = |(datain[207:204] ^ 9);
  assign w21[27] = |(datain[203:200] ^ 6);
  assign w21[28] = |(datain[199:196] ^ 14);
  assign w21[29] = |(datain[195:192] ^ 11);
  assign w21[30] = |(datain[191:188] ^ 0);
  assign w21[31] = |(datain[187:184] ^ 4);
  assign w21[32] = |(datain[183:180] ^ 12);
  assign w21[33] = |(datain[179:176] ^ 13);
  assign w21[34] = |(datain[175:172] ^ 2);
  assign w21[35] = |(datain[171:168] ^ 1);
  assign w21[36] = |(datain[167:164] ^ 5);
  assign w21[37] = |(datain[163:160] ^ 10);
  assign w21[38] = |(datain[159:156] ^ 5);
  assign w21[39] = |(datain[155:152] ^ 9);
  assign w21[40] = |(datain[151:148] ^ 8);
  assign w21[41] = |(datain[147:144] ^ 0);
  assign w21[42] = |(datain[143:140] ^ 14);
  assign w21[43] = |(datain[139:136] ^ 1);
  assign w21[44] = |(datain[135:132] ^ 14);
  assign w21[45] = |(datain[131:128] ^ 0);
  assign w21[46] = |(datain[127:124] ^ 8);
  assign w21[47] = |(datain[123:120] ^ 0);
  assign w21[48] = |(datain[119:116] ^ 12);
  assign w21[49] = |(datain[115:112] ^ 9);
  assign w21[50] = |(datain[111:108] ^ 1);
  assign w21[51] = |(datain[107:104] ^ 15);
  assign w21[52] = |(datain[103:100] ^ 11);
  assign w21[53] = |(datain[99:96] ^ 8);
  assign w21[54] = |(datain[95:92] ^ 0);
  assign w21[55] = |(datain[91:88] ^ 1);
  assign w21[56] = |(datain[87:84] ^ 5);
  assign w21[57] = |(datain[83:80] ^ 7);
  assign w21[58] = |(datain[79:76] ^ 12);
  assign w21[59] = |(datain[75:72] ^ 13);
  assign w21[60] = |(datain[71:68] ^ 2);
  assign w21[61] = |(datain[67:64] ^ 1);
  assign w21[62] = |(datain[63:60] ^ 1);
  assign w21[63] = |(datain[59:56] ^ 15);
  assign w21[64] = |(datain[55:52] ^ 5);
  assign w21[65] = |(datain[51:48] ^ 10);
  assign w21[66] = |(datain[47:44] ^ 5);
  assign w21[67] = |(datain[43:40] ^ 9);
  assign w21[68] = |(datain[39:36] ^ 14);
  assign w21[69] = |(datain[35:32] ^ 8);
  assign w21[70] = |(datain[31:28] ^ 0);
  assign w21[71] = |(datain[27:24] ^ 6);
  assign w21[72] = |(datain[23:20] ^ 0);
  assign w21[73] = |(datain[19:16] ^ 0);
  assign w21[74] = |(datain[15:12] ^ 11);
  assign w21[75] = |(datain[11:8] ^ 4);
  assign comp[21] = ~(|w21);
  wire [74-1:0] w22;
  assign w22[0] = |(datain[311:308] ^ 0);
  assign w22[1] = |(datain[307:304] ^ 14);
  assign w22[2] = |(datain[303:300] ^ 0);
  assign w22[3] = |(datain[299:296] ^ 7);
  assign w22[4] = |(datain[295:292] ^ 11);
  assign w22[5] = |(datain[291:288] ^ 9);
  assign w22[6] = |(datain[287:284] ^ 1);
  assign w22[7] = |(datain[283:280] ^ 1);
  assign w22[8] = |(datain[279:276] ^ 0);
  assign w22[9] = |(datain[275:272] ^ 0);
  assign w22[10] = |(datain[271:268] ^ 15);
  assign w22[11] = |(datain[267:264] ^ 3);
  assign w22[12] = |(datain[263:260] ^ 10);
  assign w22[13] = |(datain[259:256] ^ 4);
  assign w22[14] = |(datain[255:252] ^ 11);
  assign w22[15] = |(datain[251:248] ^ 14);
  assign w22[16] = |(datain[247:244] ^ 2);
  assign w22[17] = |(datain[243:240] ^ 14);
  assign w22[18] = |(datain[239:236] ^ 0);
  assign w22[19] = |(datain[235:232] ^ 1);
  assign w22[20] = |(datain[231:228] ^ 11);
  assign w22[21] = |(datain[227:224] ^ 9);
  assign w22[22] = |(datain[223:220] ^ 1);
  assign w22[23] = |(datain[219:216] ^ 7);
  assign w22[24] = |(datain[215:212] ^ 2);
  assign w22[25] = |(datain[211:208] ^ 2);
  assign w22[26] = |(datain[207:204] ^ 10);
  assign w22[27] = |(datain[203:200] ^ 12);
  assign w22[28] = |(datain[199:196] ^ 3);
  assign w22[29] = |(datain[195:192] ^ 2);
  assign w22[30] = |(datain[191:188] ^ 12);
  assign w22[31] = |(datain[187:184] ^ 2);
  assign w22[32] = |(datain[183:180] ^ 15);
  assign w22[33] = |(datain[179:176] ^ 6);
  assign w22[34] = |(datain[175:172] ^ 13);
  assign w22[35] = |(datain[171:168] ^ 10);
  assign w22[36] = |(datain[167:164] ^ 10);
  assign w22[37] = |(datain[163:160] ^ 10);
  assign w22[38] = |(datain[159:156] ^ 14);
  assign w22[39] = |(datain[155:152] ^ 2);
  assign w22[40] = |(datain[151:148] ^ 15);
  assign w22[41] = |(datain[147:144] ^ 8);
  assign w22[42] = |(datain[143:140] ^ 5);
  assign w22[43] = |(datain[139:136] ^ 11);
  assign w22[44] = |(datain[135:132] ^ 5);
  assign w22[45] = |(datain[131:128] ^ 15);
  assign w22[46] = |(datain[127:124] ^ 0);
  assign w22[47] = |(datain[123:120] ^ 7);
  assign w22[48] = |(datain[119:116] ^ 11);
  assign w22[49] = |(datain[115:112] ^ 4);
  assign w22[50] = |(datain[111:108] ^ 4);
  assign w22[51] = |(datain[107:104] ^ 0);
  assign w22[52] = |(datain[103:100] ^ 11);
  assign w22[53] = |(datain[99:96] ^ 9);
  assign w22[54] = |(datain[95:92] ^ 2);
  assign w22[55] = |(datain[91:88] ^ 8);
  assign w22[56] = |(datain[87:84] ^ 2);
  assign w22[57] = |(datain[83:80] ^ 2);
  assign w22[58] = |(datain[79:76] ^ 9);
  assign w22[59] = |(datain[75:72] ^ 0);
  assign w22[60] = |(datain[71:68] ^ 11);
  assign w22[61] = |(datain[67:64] ^ 10);
  assign w22[62] = |(datain[63:60] ^ 8);
  assign w22[63] = |(datain[59:56] ^ 1);
  assign w22[64] = |(datain[55:52] ^ 2);
  assign w22[65] = |(datain[51:48] ^ 3);
  assign w22[66] = |(datain[47:44] ^ 14);
  assign w22[67] = |(datain[43:40] ^ 8);
  assign w22[68] = |(datain[39:36] ^ 0);
  assign w22[69] = |(datain[35:32] ^ 4);
  assign w22[70] = |(datain[31:28] ^ 15);
  assign w22[71] = |(datain[27:24] ^ 12);
  assign w22[72] = |(datain[23:20] ^ 12);
  assign w22[73] = |(datain[19:16] ^ 3);
  assign comp[22] = ~(|w22);
  wire [76-1:0] w23;
  assign w23[0] = |(datain[311:308] ^ 0);
  assign w23[1] = |(datain[307:304] ^ 7);
  assign w23[2] = |(datain[303:300] ^ 2);
  assign w23[3] = |(datain[299:296] ^ 4);
  assign w23[4] = |(datain[295:292] ^ 5);
  assign w23[5] = |(datain[291:288] ^ 11);
  assign w23[6] = |(datain[287:284] ^ 5);
  assign w23[7] = |(datain[283:280] ^ 3);
  assign w23[8] = |(datain[279:276] ^ 11);
  assign w23[9] = |(datain[275:272] ^ 4);
  assign w23[10] = |(datain[271:268] ^ 4);
  assign w23[11] = |(datain[267:264] ^ 0);
  assign w23[12] = |(datain[263:260] ^ 11);
  assign w23[13] = |(datain[259:256] ^ 9);
  assign w23[14] = |(datain[255:252] ^ 12);
  assign w23[15] = |(datain[251:248] ^ 4);
  assign w23[16] = |(datain[247:244] ^ 0);
  assign w23[17] = |(datain[243:240] ^ 3);
  assign w23[18] = |(datain[239:236] ^ 8);
  assign w23[19] = |(datain[235:232] ^ 13);
  assign w23[20] = |(datain[231:228] ^ 9);
  assign w23[21] = |(datain[227:224] ^ 6);
  assign w23[22] = |(datain[223:220] ^ 0);
  assign w23[23] = |(datain[219:216] ^ 3);
  assign w23[24] = |(datain[215:212] ^ 0);
  assign w23[25] = |(datain[211:208] ^ 1);
  assign w23[26] = |(datain[207:204] ^ 12);
  assign w23[27] = |(datain[203:200] ^ 13);
  assign w23[28] = |(datain[199:196] ^ 2);
  assign w23[29] = |(datain[195:192] ^ 1);
  assign w23[30] = |(datain[191:188] ^ 11);
  assign w23[31] = |(datain[187:184] ^ 0);
  assign w23[32] = |(datain[183:180] ^ 0);
  assign w23[33] = |(datain[179:176] ^ 3);
  assign w23[34] = |(datain[175:172] ^ 12);
  assign w23[35] = |(datain[171:168] ^ 15);
  assign w23[36] = |(datain[167:164] ^ 11);
  assign w23[37] = |(datain[163:160] ^ 4);
  assign w23[38] = |(datain[159:156] ^ 3);
  assign w23[39] = |(datain[155:152] ^ 13);
  assign w23[40] = |(datain[151:148] ^ 8);
  assign w23[41] = |(datain[147:144] ^ 13);
  assign w23[42] = |(datain[143:140] ^ 9);
  assign w23[43] = |(datain[139:136] ^ 6);
  assign w23[44] = |(datain[135:132] ^ 4);
  assign w23[45] = |(datain[131:128] ^ 1);
  assign w23[46] = |(datain[127:124] ^ 0);
  assign w23[47] = |(datain[123:120] ^ 5);
  assign w23[48] = |(datain[119:116] ^ 12);
  assign w23[49] = |(datain[115:112] ^ 13);
  assign w23[50] = |(datain[111:108] ^ 2);
  assign w23[51] = |(datain[107:104] ^ 1);
  assign w23[52] = |(datain[103:100] ^ 9);
  assign w23[53] = |(datain[99:96] ^ 3);
  assign w23[54] = |(datain[95:92] ^ 12);
  assign w23[55] = |(datain[91:88] ^ 3);
  assign w23[56] = |(datain[87:84] ^ 11);
  assign w23[57] = |(datain[83:80] ^ 8);
  assign w23[58] = |(datain[79:76] ^ 0);
  assign w23[59] = |(datain[75:72] ^ 1);
  assign w23[60] = |(datain[71:68] ^ 4);
  assign w23[61] = |(datain[67:64] ^ 3);
  assign w23[62] = |(datain[63:60] ^ 8);
  assign w23[63] = |(datain[59:56] ^ 13);
  assign w23[64] = |(datain[55:52] ^ 9);
  assign w23[65] = |(datain[51:48] ^ 6);
  assign w23[66] = |(datain[47:44] ^ 4);
  assign w23[67] = |(datain[43:40] ^ 1);
  assign w23[68] = |(datain[39:36] ^ 0);
  assign w23[69] = |(datain[35:32] ^ 5);
  assign w23[70] = |(datain[31:28] ^ 12);
  assign w23[71] = |(datain[27:24] ^ 13);
  assign w23[72] = |(datain[23:20] ^ 2);
  assign w23[73] = |(datain[19:16] ^ 1);
  assign w23[74] = |(datain[15:12] ^ 12);
  assign w23[75] = |(datain[11:8] ^ 3);
  assign comp[23] = ~(|w23);
  wire [74-1:0] w24;
  assign w24[0] = |(datain[311:308] ^ 0);
  assign w24[1] = |(datain[307:304] ^ 14);
  assign w24[2] = |(datain[303:300] ^ 0);
  assign w24[3] = |(datain[299:296] ^ 9);
  assign w24[4] = |(datain[295:292] ^ 0);
  assign w24[5] = |(datain[291:288] ^ 1);
  assign w24[6] = |(datain[287:284] ^ 9);
  assign w24[7] = |(datain[283:280] ^ 0);
  assign w24[8] = |(datain[279:276] ^ 11);
  assign w24[9] = |(datain[275:272] ^ 10);
  assign w24[10] = |(datain[271:268] ^ 0);
  assign w24[11] = |(datain[267:264] ^ 0);
  assign w24[12] = |(datain[263:260] ^ 0);
  assign w24[13] = |(datain[259:256] ^ 1);
  assign w24[14] = |(datain[255:252] ^ 9);
  assign w24[15] = |(datain[251:248] ^ 0);
  assign w24[16] = |(datain[247:244] ^ 11);
  assign w24[17] = |(datain[243:240] ^ 4);
  assign w24[18] = |(datain[239:236] ^ 4);
  assign w24[19] = |(datain[235:232] ^ 0);
  assign w24[20] = |(datain[231:228] ^ 9);
  assign w24[21] = |(datain[227:224] ^ 0);
  assign w24[22] = |(datain[223:220] ^ 11);
  assign w24[23] = |(datain[219:216] ^ 9);
  assign w24[24] = |(datain[215:212] ^ 0);
  assign w24[25] = |(datain[211:208] ^ 13);
  assign w24[26] = |(datain[207:204] ^ 0);
  assign w24[27] = |(datain[203:200] ^ 0);
  assign w24[28] = |(datain[199:196] ^ 9);
  assign w24[29] = |(datain[195:192] ^ 0);
  assign w24[30] = |(datain[191:188] ^ 12);
  assign w24[31] = |(datain[187:184] ^ 13);
  assign w24[32] = |(datain[183:180] ^ 2);
  assign w24[33] = |(datain[179:176] ^ 1);
  assign w24[34] = |(datain[175:172] ^ 9);
  assign w24[35] = |(datain[171:168] ^ 0);
  assign w24[36] = |(datain[167:164] ^ 11);
  assign w24[37] = |(datain[163:160] ^ 8);
  assign w24[38] = |(datain[159:156] ^ 0);
  assign w24[39] = |(datain[155:152] ^ 1);
  assign w24[40] = |(datain[151:148] ^ 5);
  assign w24[41] = |(datain[147:144] ^ 7);
  assign w24[42] = |(datain[143:140] ^ 9);
  assign w24[43] = |(datain[139:136] ^ 0);
  assign w24[44] = |(datain[135:132] ^ 8);
  assign w24[45] = |(datain[131:128] ^ 11);
  assign w24[46] = |(datain[127:124] ^ 0);
  assign w24[47] = |(datain[123:120] ^ 14);
  assign w24[48] = |(datain[119:116] ^ 0);
  assign w24[49] = |(datain[115:112] ^ 9);
  assign w24[50] = |(datain[111:108] ^ 0);
  assign w24[51] = |(datain[107:104] ^ 1);
  assign w24[52] = |(datain[103:100] ^ 9);
  assign w24[53] = |(datain[99:96] ^ 0);
  assign w24[54] = |(datain[95:92] ^ 8);
  assign w24[55] = |(datain[91:88] ^ 11);
  assign w24[56] = |(datain[87:84] ^ 1);
  assign w24[57] = |(datain[83:80] ^ 6);
  assign w24[58] = |(datain[79:76] ^ 0);
  assign w24[59] = |(datain[75:72] ^ 7);
  assign w24[60] = |(datain[71:68] ^ 0);
  assign w24[61] = |(datain[67:64] ^ 1);
  assign w24[62] = |(datain[63:60] ^ 9);
  assign w24[63] = |(datain[59:56] ^ 0);
  assign w24[64] = |(datain[55:52] ^ 12);
  assign w24[65] = |(datain[51:48] ^ 13);
  assign w24[66] = |(datain[47:44] ^ 2);
  assign w24[67] = |(datain[43:40] ^ 1);
  assign w24[68] = |(datain[39:36] ^ 9);
  assign w24[69] = |(datain[35:32] ^ 0);
  assign w24[70] = |(datain[31:28] ^ 11);
  assign w24[71] = |(datain[27:24] ^ 4);
  assign w24[72] = |(datain[23:20] ^ 3);
  assign w24[73] = |(datain[19:16] ^ 14);
  assign comp[24] = ~(|w24);
  wire [74-1:0] w25;
  assign w25[0] = |(datain[311:308] ^ 8);
  assign w25[1] = |(datain[307:304] ^ 13);
  assign w25[2] = |(datain[303:300] ^ 9);
  assign w25[3] = |(datain[299:296] ^ 6);
  assign w25[4] = |(datain[295:292] ^ 5);
  assign w25[5] = |(datain[291:288] ^ 12);
  assign w25[6] = |(datain[287:284] ^ 0);
  assign w25[7] = |(datain[283:280] ^ 5);
  assign w25[8] = |(datain[279:276] ^ 12);
  assign w25[9] = |(datain[275:272] ^ 13);
  assign w25[10] = |(datain[271:268] ^ 2);
  assign w25[11] = |(datain[267:264] ^ 1);
  assign w25[12] = |(datain[263:260] ^ 3);
  assign w25[13] = |(datain[259:256] ^ 2);
  assign w25[14] = |(datain[255:252] ^ 12);
  assign w25[15] = |(datain[251:248] ^ 0);
  assign w25[16] = |(datain[247:244] ^ 14);
  assign w25[17] = |(datain[243:240] ^ 8);
  assign w25[18] = |(datain[239:236] ^ 2);
  assign w25[19] = |(datain[235:232] ^ 14);
  assign w25[20] = |(datain[231:228] ^ 0);
  assign w25[21] = |(datain[227:224] ^ 0);
  assign w25[22] = |(datain[223:220] ^ 8);
  assign w25[23] = |(datain[219:216] ^ 13);
  assign w25[24] = |(datain[215:212] ^ 9);
  assign w25[25] = |(datain[211:208] ^ 6);
  assign w25[26] = |(datain[207:204] ^ 11);
  assign w25[27] = |(datain[203:200] ^ 12);
  assign w25[28] = |(datain[199:196] ^ 0);
  assign w25[29] = |(datain[195:192] ^ 4);
  assign w25[30] = |(datain[191:188] ^ 12);
  assign w25[31] = |(datain[187:184] ^ 13);
  assign w25[32] = |(datain[183:180] ^ 2);
  assign w25[33] = |(datain[179:176] ^ 1);
  assign w25[34] = |(datain[175:172] ^ 5);
  assign w25[35] = |(datain[171:168] ^ 10);
  assign w25[36] = |(datain[167:164] ^ 5);
  assign w25[37] = |(datain[163:160] ^ 9);
  assign w25[38] = |(datain[159:156] ^ 8);
  assign w25[39] = |(datain[155:152] ^ 0);
  assign w25[40] = |(datain[151:148] ^ 14);
  assign w25[41] = |(datain[147:144] ^ 1);
  assign w25[42] = |(datain[143:140] ^ 14);
  assign w25[43] = |(datain[139:136] ^ 0);
  assign w25[44] = |(datain[135:132] ^ 8);
  assign w25[45] = |(datain[131:128] ^ 0);
  assign w25[46] = |(datain[127:124] ^ 12);
  assign w25[47] = |(datain[123:120] ^ 9);
  assign w25[48] = |(datain[119:116] ^ 0);
  assign w25[49] = |(datain[115:112] ^ 5);
  assign w25[50] = |(datain[111:108] ^ 11);
  assign w25[51] = |(datain[107:104] ^ 8);
  assign w25[52] = |(datain[103:100] ^ 0);
  assign w25[53] = |(datain[99:96] ^ 1);
  assign w25[54] = |(datain[95:92] ^ 5);
  assign w25[55] = |(datain[91:88] ^ 7);
  assign w25[56] = |(datain[87:84] ^ 12);
  assign w25[57] = |(datain[83:80] ^ 13);
  assign w25[58] = |(datain[79:76] ^ 2);
  assign w25[59] = |(datain[75:72] ^ 1);
  assign w25[60] = |(datain[71:68] ^ 3);
  assign w25[61] = |(datain[67:64] ^ 14);
  assign w25[62] = |(datain[63:60] ^ 15);
  assign w25[63] = |(datain[59:56] ^ 14);
  assign w25[64] = |(datain[55:52] ^ 8);
  assign w25[65] = |(datain[51:48] ^ 6);
  assign w25[66] = |(datain[47:44] ^ 11);
  assign w25[67] = |(datain[43:40] ^ 15);
  assign w25[68] = |(datain[39:36] ^ 0);
  assign w25[69] = |(datain[35:32] ^ 4);
  assign w25[70] = |(datain[31:28] ^ 1);
  assign w25[71] = |(datain[27:24] ^ 15);
  assign w25[72] = |(datain[23:20] ^ 5);
  assign w25[73] = |(datain[19:16] ^ 10);
  assign comp[25] = ~(|w25);
  wire [74-1:0] w26;
  assign w26[0] = |(datain[311:308] ^ 0);
  assign w26[1] = |(datain[307:304] ^ 1);
  assign w26[2] = |(datain[303:300] ^ 11);
  assign w26[3] = |(datain[299:296] ^ 9);
  assign w26[4] = |(datain[295:292] ^ 1);
  assign w26[5] = |(datain[291:288] ^ 9);
  assign w26[6] = |(datain[287:284] ^ 0);
  assign w26[7] = |(datain[283:280] ^ 0);
  assign w26[8] = |(datain[279:276] ^ 12);
  assign w26[9] = |(datain[275:272] ^ 13);
  assign w26[10] = |(datain[271:268] ^ 2);
  assign w26[11] = |(datain[267:264] ^ 1);
  assign w26[12] = |(datain[263:260] ^ 11);
  assign w26[13] = |(datain[259:256] ^ 4);
  assign w26[14] = |(datain[255:252] ^ 4);
  assign w26[15] = |(datain[251:248] ^ 0);
  assign w26[16] = |(datain[247:244] ^ 8);
  assign w26[17] = |(datain[243:240] ^ 13);
  assign w26[18] = |(datain[239:236] ^ 9);
  assign w26[19] = |(datain[235:232] ^ 6);
  assign w26[20] = |(datain[231:228] ^ 2);
  assign w26[21] = |(datain[227:224] ^ 2);
  assign w26[22] = |(datain[223:220] ^ 0);
  assign w26[23] = |(datain[219:216] ^ 3);
  assign w26[24] = |(datain[215:212] ^ 11);
  assign w26[25] = |(datain[211:208] ^ 9);
  assign w26[26] = |(datain[207:204] ^ 15);
  assign w26[27] = |(datain[203:200] ^ 8);
  assign w26[28] = |(datain[199:196] ^ 0);
  assign w26[29] = |(datain[195:192] ^ 1);
  assign w26[30] = |(datain[191:188] ^ 12);
  assign w26[31] = |(datain[187:184] ^ 13);
  assign w26[32] = |(datain[183:180] ^ 2);
  assign w26[33] = |(datain[179:176] ^ 1);
  assign w26[34] = |(datain[175:172] ^ 11);
  assign w26[35] = |(datain[171:168] ^ 4);
  assign w26[36] = |(datain[167:164] ^ 4);
  assign w26[37] = |(datain[163:160] ^ 0);
  assign w26[38] = |(datain[159:156] ^ 8);
  assign w26[39] = |(datain[155:152] ^ 13);
  assign w26[40] = |(datain[151:148] ^ 9);
  assign w26[41] = |(datain[147:144] ^ 6);
  assign w26[42] = |(datain[143:140] ^ 1);
  assign w26[43] = |(datain[139:136] ^ 4);
  assign w26[44] = |(datain[135:132] ^ 0);
  assign w26[45] = |(datain[131:128] ^ 3);
  assign w26[46] = |(datain[127:124] ^ 11);
  assign w26[47] = |(datain[123:120] ^ 9);
  assign w26[48] = |(datain[119:116] ^ 0);
  assign w26[49] = |(datain[115:112] ^ 14);
  assign w26[50] = |(datain[111:108] ^ 0);
  assign w26[51] = |(datain[107:104] ^ 0);
  assign w26[52] = |(datain[103:100] ^ 12);
  assign w26[53] = |(datain[99:96] ^ 13);
  assign w26[54] = |(datain[95:92] ^ 2);
  assign w26[55] = |(datain[91:88] ^ 1);
  assign w26[56] = |(datain[87:84] ^ 5);
  assign w26[57] = |(datain[83:80] ^ 9);
  assign w26[58] = |(datain[79:76] ^ 8);
  assign w26[59] = |(datain[75:72] ^ 8);
  assign w26[60] = |(datain[71:68] ^ 8);
  assign w26[61] = |(datain[67:64] ^ 14);
  assign w26[62] = |(datain[63:60] ^ 1);
  assign w26[63] = |(datain[59:56] ^ 1);
  assign w26[64] = |(datain[55:52] ^ 0);
  assign w26[65] = |(datain[51:48] ^ 3);
  assign w26[66] = |(datain[47:44] ^ 8);
  assign w26[67] = |(datain[43:40] ^ 0);
  assign w26[68] = |(datain[39:36] ^ 10);
  assign w26[69] = |(datain[35:32] ^ 14);
  assign w26[70] = |(datain[31:28] ^ 1);
  assign w26[71] = |(datain[27:24] ^ 1);
  assign w26[72] = |(datain[23:20] ^ 0);
  assign w26[73] = |(datain[19:16] ^ 3);
  assign comp[26] = ~(|w26);
  wire [76-1:0] w27;
  assign w27[0] = |(datain[311:308] ^ 2);
  assign w27[1] = |(datain[307:304] ^ 2);
  assign w27[2] = |(datain[303:300] ^ 0);
  assign w27[3] = |(datain[299:296] ^ 3);
  assign w27[4] = |(datain[295:292] ^ 11);
  assign w27[5] = |(datain[291:288] ^ 9);
  assign w27[6] = |(datain[287:284] ^ 15);
  assign w27[7] = |(datain[283:280] ^ 8);
  assign w27[8] = |(datain[279:276] ^ 0);
  assign w27[9] = |(datain[275:272] ^ 1);
  assign w27[10] = |(datain[271:268] ^ 12);
  assign w27[11] = |(datain[267:264] ^ 13);
  assign w27[12] = |(datain[263:260] ^ 2);
  assign w27[13] = |(datain[259:256] ^ 1);
  assign w27[14] = |(datain[255:252] ^ 11);
  assign w27[15] = |(datain[251:248] ^ 4);
  assign w27[16] = |(datain[247:244] ^ 4);
  assign w27[17] = |(datain[243:240] ^ 0);
  assign w27[18] = |(datain[239:236] ^ 8);
  assign w27[19] = |(datain[235:232] ^ 13);
  assign w27[20] = |(datain[231:228] ^ 9);
  assign w27[21] = |(datain[227:224] ^ 6);
  assign w27[22] = |(datain[223:220] ^ 1);
  assign w27[23] = |(datain[219:216] ^ 4);
  assign w27[24] = |(datain[215:212] ^ 0);
  assign w27[25] = |(datain[211:208] ^ 3);
  assign w27[26] = |(datain[207:204] ^ 11);
  assign w27[27] = |(datain[203:200] ^ 9);
  assign w27[28] = |(datain[199:196] ^ 0);
  assign w27[29] = |(datain[195:192] ^ 14);
  assign w27[30] = |(datain[191:188] ^ 0);
  assign w27[31] = |(datain[187:184] ^ 0);
  assign w27[32] = |(datain[183:180] ^ 12);
  assign w27[33] = |(datain[179:176] ^ 13);
  assign w27[34] = |(datain[175:172] ^ 2);
  assign w27[35] = |(datain[171:168] ^ 1);
  assign w27[36] = |(datain[167:164] ^ 5);
  assign w27[37] = |(datain[163:160] ^ 9);
  assign w27[38] = |(datain[159:156] ^ 8);
  assign w27[39] = |(datain[155:152] ^ 8);
  assign w27[40] = |(datain[151:148] ^ 8);
  assign w27[41] = |(datain[147:144] ^ 14);
  assign w27[42] = |(datain[143:140] ^ 1);
  assign w27[43] = |(datain[139:136] ^ 1);
  assign w27[44] = |(datain[135:132] ^ 0);
  assign w27[45] = |(datain[131:128] ^ 3);
  assign w27[46] = |(datain[127:124] ^ 8);
  assign w27[47] = |(datain[123:120] ^ 0);
  assign w27[48] = |(datain[119:116] ^ 10);
  assign w27[49] = |(datain[115:112] ^ 14);
  assign w27[50] = |(datain[111:108] ^ 1);
  assign w27[51] = |(datain[107:104] ^ 1);
  assign w27[52] = |(datain[103:100] ^ 0);
  assign w27[53] = |(datain[99:96] ^ 3);
  assign w27[54] = |(datain[95:92] ^ 0);
  assign w27[55] = |(datain[91:88] ^ 1);
  assign w27[56] = |(datain[87:84] ^ 8);
  assign w27[57] = |(datain[83:80] ^ 0);
  assign w27[58] = |(datain[79:76] ^ 11);
  assign w27[59] = |(datain[75:72] ^ 14);
  assign w27[60] = |(datain[71:68] ^ 1);
  assign w27[61] = |(datain[67:64] ^ 1);
  assign w27[62] = |(datain[63:60] ^ 0);
  assign w27[63] = |(datain[59:56] ^ 3);
  assign w27[64] = |(datain[55:52] ^ 0);
  assign w27[65] = |(datain[51:48] ^ 0);
  assign w27[66] = |(datain[47:44] ^ 7);
  assign w27[67] = |(datain[43:40] ^ 4);
  assign w27[68] = |(datain[39:36] ^ 2);
  assign w27[69] = |(datain[35:32] ^ 3);
  assign w27[70] = |(datain[31:28] ^ 11);
  assign w27[71] = |(datain[27:24] ^ 8);
  assign w27[72] = |(datain[23:20] ^ 0);
  assign w27[73] = |(datain[19:16] ^ 1);
  assign w27[74] = |(datain[15:12] ^ 5);
  assign w27[75] = |(datain[11:8] ^ 7);
  assign comp[27] = ~(|w27);
  wire [76-1:0] w28;
  assign w28[0] = |(datain[311:308] ^ 15);
  assign w28[1] = |(datain[307:304] ^ 10);
  assign w28[2] = |(datain[303:300] ^ 2);
  assign w28[3] = |(datain[299:296] ^ 6);
  assign w28[4] = |(datain[295:292] ^ 10);
  assign w28[5] = |(datain[291:288] ^ 3);
  assign w28[6] = |(datain[287:284] ^ 9);
  assign w28[7] = |(datain[283:280] ^ 0);
  assign w28[8] = |(datain[279:276] ^ 0);
  assign w28[9] = |(datain[275:272] ^ 0);
  assign w28[10] = |(datain[271:268] ^ 2);
  assign w28[11] = |(datain[267:264] ^ 6);
  assign w28[12] = |(datain[263:260] ^ 8);
  assign w28[13] = |(datain[259:256] ^ 9);
  assign w28[14] = |(datain[255:252] ^ 1);
  assign w28[15] = |(datain[251:248] ^ 14);
  assign w28[16] = |(datain[247:244] ^ 9);
  assign w28[17] = |(datain[243:240] ^ 2);
  assign w28[18] = |(datain[239:236] ^ 0);
  assign w28[19] = |(datain[235:232] ^ 0);
  assign w28[20] = |(datain[231:228] ^ 15);
  assign w28[21] = |(datain[227:224] ^ 11);
  assign w28[22] = |(datain[223:220] ^ 12);
  assign w28[23] = |(datain[219:216] ^ 3);
  assign w28[24] = |(datain[215:212] ^ 9);
  assign w28[25] = |(datain[211:208] ^ 12);
  assign w28[26] = |(datain[207:204] ^ 2);
  assign w28[27] = |(datain[203:200] ^ 14);
  assign w28[28] = |(datain[199:196] ^ 15);
  assign w28[29] = |(datain[195:192] ^ 15);
  assign w28[30] = |(datain[191:188] ^ 1);
  assign w28[31] = |(datain[187:184] ^ 14);
  assign w28[32] = |(datain[183:180] ^ 0);
  assign w28[33] = |(datain[179:176] ^ 2);
  assign w28[34] = |(datain[175:172] ^ 0);
  assign w28[35] = |(datain[171:168] ^ 5);
  assign w28[36] = |(datain[167:164] ^ 12);
  assign w28[37] = |(datain[163:160] ^ 3);
  assign w28[38] = |(datain[159:156] ^ 11);
  assign w28[39] = |(datain[155:152] ^ 8);
  assign w28[40] = |(datain[151:148] ^ 0);
  assign w28[41] = |(datain[147:144] ^ 0);
  assign w28[42] = |(datain[143:140] ^ 4);
  assign w28[43] = |(datain[139:136] ^ 2);
  assign w28[44] = |(datain[135:132] ^ 3);
  assign w28[45] = |(datain[131:128] ^ 3);
  assign w28[46] = |(datain[127:124] ^ 12);
  assign w28[47] = |(datain[123:120] ^ 9);
  assign w28[48] = |(datain[119:116] ^ 3);
  assign w28[49] = |(datain[115:112] ^ 3);
  assign w28[50] = |(datain[111:108] ^ 13);
  assign w28[51] = |(datain[107:104] ^ 2);
  assign w28[52] = |(datain[103:100] ^ 14);
  assign w28[53] = |(datain[99:96] ^ 8);
  assign w28[54] = |(datain[95:92] ^ 14);
  assign w28[55] = |(datain[91:88] ^ 15);
  assign w28[56] = |(datain[87:84] ^ 15);
  assign w28[57] = |(datain[83:80] ^ 15);
  assign w28[58] = |(datain[79:76] ^ 12);
  assign w28[59] = |(datain[75:72] ^ 3);
  assign w28[60] = |(datain[71:68] ^ 11);
  assign w28[61] = |(datain[67:64] ^ 4);
  assign w28[62] = |(datain[63:60] ^ 3);
  assign w28[63] = |(datain[59:56] ^ 14);
  assign w28[64] = |(datain[55:52] ^ 14);
  assign w28[65] = |(datain[51:48] ^ 8);
  assign w28[66] = |(datain[47:44] ^ 14);
  assign w28[67] = |(datain[43:40] ^ 9);
  assign w28[68] = |(datain[39:36] ^ 15);
  assign w28[69] = |(datain[35:32] ^ 15);
  assign w28[70] = |(datain[31:28] ^ 12);
  assign w28[71] = |(datain[27:24] ^ 3);
  assign w28[72] = |(datain[23:20] ^ 10);
  assign w28[73] = |(datain[19:16] ^ 1);
  assign w28[74] = |(datain[15:12] ^ 1);
  assign w28[75] = |(datain[11:8] ^ 13);
  assign comp[28] = ~(|w28);
  wire [76-1:0] w29;
  assign w29[0] = |(datain[311:308] ^ 12);
  assign w29[1] = |(datain[307:304] ^ 13);
  assign w29[2] = |(datain[303:300] ^ 2);
  assign w29[3] = |(datain[299:296] ^ 1);
  assign w29[4] = |(datain[295:292] ^ 11);
  assign w29[5] = |(datain[291:288] ^ 10);
  assign w29[6] = |(datain[287:284] ^ 9);
  assign w29[7] = |(datain[283:280] ^ 3);
  assign w29[8] = |(datain[279:276] ^ 0);
  assign w29[9] = |(datain[275:272] ^ 5);
  assign w29[10] = |(datain[271:268] ^ 11);
  assign w29[11] = |(datain[267:264] ^ 13);
  assign w29[12] = |(datain[263:260] ^ 0);
  assign w29[13] = |(datain[259:256] ^ 10);
  assign w29[14] = |(datain[255:252] ^ 0);
  assign w29[15] = |(datain[251:248] ^ 0);
  assign w29[16] = |(datain[247:244] ^ 3);
  assign w29[17] = |(datain[243:240] ^ 3);
  assign w29[18] = |(datain[239:236] ^ 12);
  assign w29[19] = |(datain[235:232] ^ 9);
  assign w29[20] = |(datain[231:228] ^ 11);
  assign w29[21] = |(datain[227:224] ^ 4);
  assign w29[22] = |(datain[223:220] ^ 3);
  assign w29[23] = |(datain[219:216] ^ 12);
  assign w29[24] = |(datain[215:212] ^ 12);
  assign w29[25] = |(datain[211:208] ^ 13);
  assign w29[26] = |(datain[207:204] ^ 2);
  assign w29[27] = |(datain[203:200] ^ 1);
  assign w29[28] = |(datain[199:196] ^ 7);
  assign w29[29] = |(datain[195:192] ^ 2);
  assign w29[30] = |(datain[191:188] ^ 0);
  assign w29[31] = |(datain[187:184] ^ 5);
  assign w29[32] = |(datain[183:180] ^ 9);
  assign w29[33] = |(datain[179:176] ^ 3);
  assign w29[34] = |(datain[175:172] ^ 11);
  assign w29[35] = |(datain[171:168] ^ 4);
  assign w29[36] = |(datain[167:164] ^ 3);
  assign w29[37] = |(datain[163:160] ^ 14);
  assign w29[38] = |(datain[159:156] ^ 12);
  assign w29[39] = |(datain[155:152] ^ 13);
  assign w29[40] = |(datain[151:148] ^ 2);
  assign w29[41] = |(datain[147:144] ^ 1);
  assign w29[42] = |(datain[143:140] ^ 8);
  assign w29[43] = |(datain[139:136] ^ 3);
  assign w29[44] = |(datain[135:132] ^ 12);
  assign w29[45] = |(datain[131:128] ^ 2);
  assign w29[46] = |(datain[127:124] ^ 0);
  assign w29[47] = |(datain[123:120] ^ 9);
  assign w29[48] = |(datain[119:116] ^ 4);
  assign w29[49] = |(datain[115:112] ^ 13);
  assign w29[50] = |(datain[111:108] ^ 7);
  assign w29[51] = |(datain[107:104] ^ 5);
  assign w29[52] = |(datain[103:100] ^ 14);
  assign w29[53] = |(datain[99:96] ^ 13);
  assign w29[54] = |(datain[95:92] ^ 11);
  assign w29[55] = |(datain[91:88] ^ 10);
  assign w29[56] = |(datain[87:84] ^ 9);
  assign w29[57] = |(datain[83:80] ^ 0);
  assign w29[58] = |(datain[79:76] ^ 0);
  assign w29[59] = |(datain[75:72] ^ 5);
  assign w29[60] = |(datain[71:68] ^ 11);
  assign w29[61] = |(datain[67:64] ^ 4);
  assign w29[62] = |(datain[63:60] ^ 3);
  assign w29[63] = |(datain[59:56] ^ 11);
  assign w29[64] = |(datain[55:52] ^ 12);
  assign w29[65] = |(datain[51:48] ^ 13);
  assign w29[66] = |(datain[47:44] ^ 2);
  assign w29[67] = |(datain[43:40] ^ 1);
  assign w29[68] = |(datain[39:36] ^ 8);
  assign w29[69] = |(datain[35:32] ^ 0);
  assign w29[70] = |(datain[31:28] ^ 3);
  assign w29[71] = |(datain[27:24] ^ 14);
  assign w29[72] = |(datain[23:20] ^ 1);
  assign w29[73] = |(datain[19:16] ^ 1);
  assign w29[74] = |(datain[15:12] ^ 0);
  assign w29[75] = |(datain[11:8] ^ 7);
  assign comp[29] = ~(|w29);
  wire [74-1:0] w30;
  assign w30[0] = |(datain[311:308] ^ 3);
  assign w30[1] = |(datain[307:304] ^ 3);
  assign w30[2] = |(datain[303:300] ^ 12);
  assign w30[3] = |(datain[299:296] ^ 9);
  assign w30[4] = |(datain[295:292] ^ 3);
  assign w30[5] = |(datain[291:288] ^ 3);
  assign w30[6] = |(datain[287:284] ^ 13);
  assign w30[7] = |(datain[283:280] ^ 2);
  assign w30[8] = |(datain[279:276] ^ 12);
  assign w30[9] = |(datain[275:272] ^ 13);
  assign w30[10] = |(datain[271:268] ^ 2);
  assign w30[11] = |(datain[267:264] ^ 1);
  assign w30[12] = |(datain[263:260] ^ 10);
  assign w30[13] = |(datain[259:256] ^ 1);
  assign w30[14] = |(datain[255:252] ^ 2);
  assign w30[15] = |(datain[251:248] ^ 8);
  assign w30[16] = |(datain[247:244] ^ 0);
  assign w30[17] = |(datain[243:240] ^ 6);
  assign w30[18] = |(datain[239:236] ^ 2);
  assign w30[19] = |(datain[235:232] ^ 13);
  assign w30[20] = |(datain[231:228] ^ 0);
  assign w30[21] = |(datain[227:224] ^ 5);
  assign w30[22] = |(datain[223:220] ^ 0);
  assign w30[23] = |(datain[219:216] ^ 0);
  assign w30[24] = |(datain[215:212] ^ 10);
  assign w30[25] = |(datain[211:208] ^ 3);
  assign w30[26] = |(datain[207:204] ^ 2);
  assign w30[27] = |(datain[203:200] ^ 13);
  assign w30[28] = |(datain[199:196] ^ 0);
  assign w30[29] = |(datain[195:192] ^ 1);
  assign w30[30] = |(datain[191:188] ^ 11);
  assign w30[31] = |(datain[187:184] ^ 4);
  assign w30[32] = |(datain[183:180] ^ 4);
  assign w30[33] = |(datain[179:176] ^ 0);
  assign w30[34] = |(datain[175:172] ^ 11);
  assign w30[35] = |(datain[171:168] ^ 9);
  assign w30[36] = |(datain[167:164] ^ 0);
  assign w30[37] = |(datain[163:160] ^ 6);
  assign w30[38] = |(datain[159:156] ^ 0);
  assign w30[39] = |(datain[155:152] ^ 0);
  assign w30[40] = |(datain[151:148] ^ 11);
  assign w30[41] = |(datain[147:144] ^ 10);
  assign w30[42] = |(datain[143:140] ^ 2);
  assign w30[43] = |(datain[139:136] ^ 10);
  assign w30[44] = |(datain[135:132] ^ 0);
  assign w30[45] = |(datain[131:128] ^ 1);
  assign w30[46] = |(datain[127:124] ^ 12);
  assign w30[47] = |(datain[123:120] ^ 13);
  assign w30[48] = |(datain[119:116] ^ 2);
  assign w30[49] = |(datain[115:112] ^ 1);
  assign w30[50] = |(datain[111:108] ^ 11);
  assign w30[51] = |(datain[107:104] ^ 8);
  assign w30[52] = |(datain[103:100] ^ 0);
  assign w30[53] = |(datain[99:96] ^ 2);
  assign w30[54] = |(datain[95:92] ^ 4);
  assign w30[55] = |(datain[91:88] ^ 2);
  assign w30[56] = |(datain[87:84] ^ 3);
  assign w30[57] = |(datain[83:80] ^ 3);
  assign w30[58] = |(datain[79:76] ^ 12);
  assign w30[59] = |(datain[75:72] ^ 9);
  assign w30[60] = |(datain[71:68] ^ 3);
  assign w30[61] = |(datain[67:64] ^ 3);
  assign w30[62] = |(datain[63:60] ^ 13);
  assign w30[63] = |(datain[59:56] ^ 2);
  assign w30[64] = |(datain[55:52] ^ 12);
  assign w30[65] = |(datain[51:48] ^ 13);
  assign w30[66] = |(datain[47:44] ^ 2);
  assign w30[67] = |(datain[43:40] ^ 1);
  assign w30[68] = |(datain[39:36] ^ 5);
  assign w30[69] = |(datain[35:32] ^ 3);
  assign w30[70] = |(datain[31:28] ^ 10);
  assign w30[71] = |(datain[27:24] ^ 1);
  assign w30[72] = |(datain[23:20] ^ 0);
  assign w30[73] = |(datain[19:16] ^ 7);
  assign comp[30] = ~(|w30);
  wire [76-1:0] w31;
  assign w31[0] = |(datain[311:308] ^ 0);
  assign w31[1] = |(datain[307:304] ^ 3);
  assign w31[2] = |(datain[303:300] ^ 0);
  assign w31[3] = |(datain[299:296] ^ 1);
  assign w31[4] = |(datain[295:292] ^ 8);
  assign w31[5] = |(datain[291:288] ^ 9);
  assign w31[6] = |(datain[287:284] ^ 1);
  assign w31[7] = |(datain[283:280] ^ 6);
  assign w31[8] = |(datain[279:276] ^ 1);
  assign w31[9] = |(datain[275:272] ^ 9);
  assign w31[10] = |(datain[271:268] ^ 0);
  assign w31[11] = |(datain[267:264] ^ 4);
  assign w31[12] = |(datain[263:260] ^ 0);
  assign w31[13] = |(datain[259:256] ^ 14);
  assign w31[14] = |(datain[255:252] ^ 0);
  assign w31[15] = |(datain[251:248] ^ 7);
  assign w31[16] = |(datain[247:244] ^ 11);
  assign w31[17] = |(datain[243:240] ^ 9);
  assign w31[18] = |(datain[239:236] ^ 1);
  assign w31[19] = |(datain[235:232] ^ 8);
  assign w31[20] = |(datain[231:228] ^ 0);
  assign w31[21] = |(datain[227:224] ^ 4);
  assign w31[22] = |(datain[223:220] ^ 11);
  assign w31[23] = |(datain[219:216] ^ 15);
  assign w31[24] = |(datain[215:212] ^ 3);
  assign w31[25] = |(datain[211:208] ^ 10);
  assign w31[26] = |(datain[207:204] ^ 0);
  assign w31[27] = |(datain[203:200] ^ 4);
  assign w31[28] = |(datain[199:196] ^ 11);
  assign w31[29] = |(datain[195:192] ^ 14);
  assign w31[30] = |(datain[191:188] ^ 0);
  assign w31[31] = |(datain[187:184] ^ 6);
  assign w31[32] = |(datain[183:180] ^ 0);
  assign w31[33] = |(datain[179:176] ^ 0);
  assign w31[34] = |(datain[175:172] ^ 14);
  assign w31[35] = |(datain[171:168] ^ 8);
  assign w31[36] = |(datain[167:164] ^ 10);
  assign w31[37] = |(datain[163:160] ^ 9);
  assign w31[38] = |(datain[159:156] ^ 0);
  assign w31[39] = |(datain[155:152] ^ 0);
  assign w31[40] = |(datain[151:148] ^ 5);
  assign w31[41] = |(datain[147:144] ^ 1);
  assign w31[42] = |(datain[143:140] ^ 11);
  assign w31[43] = |(datain[139:136] ^ 9);
  assign w31[44] = |(datain[135:132] ^ 0);
  assign w31[45] = |(datain[131:128] ^ 3);
  assign w31[46] = |(datain[127:124] ^ 0);
  assign w31[47] = |(datain[123:120] ^ 0);
  assign w31[48] = |(datain[119:116] ^ 11);
  assign w31[49] = |(datain[115:112] ^ 4);
  assign w31[50] = |(datain[111:108] ^ 4);
  assign w31[51] = |(datain[107:104] ^ 0);
  assign w31[52] = |(datain[103:100] ^ 11);
  assign w31[53] = |(datain[99:96] ^ 10);
  assign w31[54] = |(datain[95:92] ^ 1);
  assign w31[55] = |(datain[91:88] ^ 14);
  assign w31[56] = |(datain[87:84] ^ 0);
  assign w31[57] = |(datain[83:80] ^ 4);
  assign w31[58] = |(datain[79:76] ^ 12);
  assign w31[59] = |(datain[75:72] ^ 13);
  assign w31[60] = |(datain[71:68] ^ 2);
  assign w31[61] = |(datain[67:64] ^ 1);
  assign w31[62] = |(datain[63:60] ^ 11);
  assign w31[63] = |(datain[59:56] ^ 4);
  assign w31[64] = |(datain[55:52] ^ 4);
  assign w31[65] = |(datain[51:48] ^ 0);
  assign w31[66] = |(datain[47:44] ^ 5);
  assign w31[67] = |(datain[43:40] ^ 9);
  assign w31[68] = |(datain[39:36] ^ 11);
  assign w31[69] = |(datain[35:32] ^ 10);
  assign w31[70] = |(datain[31:28] ^ 3);
  assign w31[71] = |(datain[27:24] ^ 10);
  assign w31[72] = |(datain[23:20] ^ 0);
  assign w31[73] = |(datain[19:16] ^ 4);
  assign w31[74] = |(datain[15:12] ^ 12);
  assign w31[75] = |(datain[11:8] ^ 13);
  assign comp[31] = ~(|w31);
  wire [74-1:0] w32;
  assign w32[0] = |(datain[311:308] ^ 11);
  assign w32[1] = |(datain[307:304] ^ 10);
  assign w32[2] = |(datain[303:300] ^ 8);
  assign w32[3] = |(datain[299:296] ^ 5);
  assign w32[4] = |(datain[295:292] ^ 0);
  assign w32[5] = |(datain[291:288] ^ 14);
  assign w32[6] = |(datain[287:284] ^ 11);
  assign w32[7] = |(datain[283:280] ^ 4);
  assign w32[8] = |(datain[279:276] ^ 4);
  assign w32[9] = |(datain[275:272] ^ 0);
  assign w32[10] = |(datain[271:268] ^ 14);
  assign w32[11] = |(datain[267:264] ^ 8);
  assign w32[12] = |(datain[263:260] ^ 9);
  assign w32[13] = |(datain[259:256] ^ 2);
  assign w32[14] = |(datain[255:252] ^ 0);
  assign w32[15] = |(datain[251:248] ^ 4);
  assign w32[16] = |(datain[247:244] ^ 7);
  assign w32[17] = |(datain[243:240] ^ 2);
  assign w32[18] = |(datain[239:236] ^ 1);
  assign w32[19] = |(datain[235:232] ^ 12);
  assign w32[20] = |(datain[231:228] ^ 11);
  assign w32[21] = |(datain[227:224] ^ 10);
  assign w32[22] = |(datain[223:220] ^ 7);
  assign w32[23] = |(datain[219:216] ^ 13);
  assign w32[24] = |(datain[215:212] ^ 0);
  assign w32[25] = |(datain[211:208] ^ 13);
  assign w32[26] = |(datain[207:204] ^ 11);
  assign w32[27] = |(datain[203:200] ^ 9);
  assign w32[28] = |(datain[199:196] ^ 1);
  assign w32[29] = |(datain[195:192] ^ 12);
  assign w32[30] = |(datain[191:188] ^ 0);
  assign w32[31] = |(datain[187:184] ^ 0);
  assign w32[32] = |(datain[183:180] ^ 11);
  assign w32[33] = |(datain[179:176] ^ 4);
  assign w32[34] = |(datain[175:172] ^ 4);
  assign w32[35] = |(datain[171:168] ^ 0);
  assign w32[36] = |(datain[167:164] ^ 14);
  assign w32[37] = |(datain[163:160] ^ 8);
  assign w32[38] = |(datain[159:156] ^ 8);
  assign w32[39] = |(datain[155:152] ^ 5);
  assign w32[40] = |(datain[151:148] ^ 0);
  assign w32[41] = |(datain[147:144] ^ 4);
  assign w32[42] = |(datain[143:140] ^ 14);
  assign w32[43] = |(datain[139:136] ^ 8);
  assign w32[44] = |(datain[135:132] ^ 14);
  assign w32[45] = |(datain[131:128] ^ 6);
  assign w32[46] = |(datain[127:124] ^ 0);
  assign w32[47] = |(datain[123:120] ^ 0);
  assign w32[48] = |(datain[119:116] ^ 11);
  assign w32[49] = |(datain[115:112] ^ 10);
  assign w32[50] = |(datain[111:108] ^ 7);
  assign w32[51] = |(datain[107:104] ^ 10);
  assign w32[52] = |(datain[103:100] ^ 0);
  assign w32[53] = |(datain[99:96] ^ 13);
  assign w32[54] = |(datain[95:92] ^ 11);
  assign w32[55] = |(datain[91:88] ^ 9);
  assign w32[56] = |(datain[87:84] ^ 0);
  assign w32[57] = |(datain[83:80] ^ 3);
  assign w32[58] = |(datain[79:76] ^ 0);
  assign w32[59] = |(datain[75:72] ^ 0);
  assign w32[60] = |(datain[71:68] ^ 11);
  assign w32[61] = |(datain[67:64] ^ 4);
  assign w32[62] = |(datain[63:60] ^ 4);
  assign w32[63] = |(datain[59:56] ^ 0);
  assign w32[64] = |(datain[55:52] ^ 14);
  assign w32[65] = |(datain[51:48] ^ 8);
  assign w32[66] = |(datain[47:44] ^ 7);
  assign w32[67] = |(datain[43:40] ^ 7);
  assign w32[68] = |(datain[39:36] ^ 0);
  assign w32[69] = |(datain[35:32] ^ 4);
  assign w32[70] = |(datain[31:28] ^ 14);
  assign w32[71] = |(datain[27:24] ^ 8);
  assign w32[72] = |(datain[23:20] ^ 1);
  assign w32[73] = |(datain[19:16] ^ 14);
  assign comp[32] = ~(|w32);
  wire [76-1:0] w33;
  assign w33[0] = |(datain[311:308] ^ 10);
  assign w33[1] = |(datain[307:304] ^ 2);
  assign w33[2] = |(datain[303:300] ^ 0);
  assign w33[3] = |(datain[299:296] ^ 9);
  assign w33[4] = |(datain[295:292] ^ 8);
  assign w33[5] = |(datain[291:288] ^ 11);
  assign w33[6] = |(datain[287:284] ^ 13);
  assign w33[7] = |(datain[283:280] ^ 0);
  assign w33[8] = |(datain[279:276] ^ 8);
  assign w33[9] = |(datain[275:272] ^ 1);
  assign w33[10] = |(datain[271:268] ^ 12);
  assign w33[11] = |(datain[267:264] ^ 2);
  assign w33[12] = |(datain[263:260] ^ 0);
  assign w33[13] = |(datain[259:256] ^ 0);
  assign w33[14] = |(datain[255:252] ^ 0);
  assign w33[15] = |(datain[251:248] ^ 1);
  assign w33[16] = |(datain[247:244] ^ 11);
  assign w33[17] = |(datain[243:240] ^ 0);
  assign w33[18] = |(datain[239:236] ^ 0);
  assign w33[19] = |(datain[235:232] ^ 7);
  assign w33[20] = |(datain[231:228] ^ 14);
  assign w33[21] = |(datain[227:224] ^ 8);
  assign w33[22] = |(datain[223:220] ^ 11);
  assign w33[23] = |(datain[219:216] ^ 1);
  assign w33[24] = |(datain[215:212] ^ 0);
  assign w33[25] = |(datain[211:208] ^ 1);
  assign w33[26] = |(datain[207:204] ^ 5);
  assign w33[27] = |(datain[203:200] ^ 10);
  assign w33[28] = |(datain[199:196] ^ 11);
  assign w33[29] = |(datain[195:192] ^ 4);
  assign w33[30] = |(datain[191:188] ^ 4);
  assign w33[31] = |(datain[187:184] ^ 0);
  assign w33[32] = |(datain[183:180] ^ 12);
  assign w33[33] = |(datain[179:176] ^ 13);
  assign w33[34] = |(datain[175:172] ^ 2);
  assign w33[35] = |(datain[171:168] ^ 1);
  assign w33[36] = |(datain[167:164] ^ 14);
  assign w33[37] = |(datain[163:160] ^ 8);
  assign w33[38] = |(datain[159:156] ^ 12);
  assign w33[39] = |(datain[155:152] ^ 6);
  assign w33[40] = |(datain[151:148] ^ 0);
  assign w33[41] = |(datain[147:144] ^ 0);
  assign w33[42] = |(datain[143:140] ^ 5);
  assign w33[43] = |(datain[139:136] ^ 8);
  assign w33[44] = |(datain[135:132] ^ 2);
  assign w33[45] = |(datain[131:128] ^ 13);
  assign w33[46] = |(datain[127:124] ^ 0);
  assign w33[47] = |(datain[123:120] ^ 3);
  assign w33[48] = |(datain[119:116] ^ 0);
  assign w33[49] = |(datain[115:112] ^ 0);
  assign w33[50] = |(datain[111:108] ^ 10);
  assign w33[51] = |(datain[107:104] ^ 3);
  assign w33[52] = |(datain[103:100] ^ 10);
  assign w33[53] = |(datain[99:96] ^ 2);
  assign w33[54] = |(datain[95:92] ^ 0);
  assign w33[55] = |(datain[91:88] ^ 2);
  assign w33[56] = |(datain[87:84] ^ 11);
  assign w33[57] = |(datain[83:80] ^ 10);
  assign w33[58] = |(datain[79:76] ^ 10);
  assign w33[59] = |(datain[75:72] ^ 1);
  assign w33[60] = |(datain[71:68] ^ 0);
  assign w33[61] = |(datain[67:64] ^ 2);
  assign w33[62] = |(datain[63:60] ^ 11);
  assign w33[63] = |(datain[59:56] ^ 9);
  assign w33[64] = |(datain[55:52] ^ 0);
  assign w33[65] = |(datain[51:48] ^ 4);
  assign w33[66] = |(datain[47:44] ^ 0);
  assign w33[67] = |(datain[43:40] ^ 0);
  assign w33[68] = |(datain[39:36] ^ 11);
  assign w33[69] = |(datain[35:32] ^ 4);
  assign w33[70] = |(datain[31:28] ^ 4);
  assign w33[71] = |(datain[27:24] ^ 0);
  assign w33[72] = |(datain[23:20] ^ 12);
  assign w33[73] = |(datain[19:16] ^ 13);
  assign w33[74] = |(datain[15:12] ^ 2);
  assign w33[75] = |(datain[11:8] ^ 1);
  assign comp[33] = ~(|w33);
  wire [74-1:0] w34;
  assign w34[0] = |(datain[311:308] ^ 12);
  assign w34[1] = |(datain[307:304] ^ 1);
  assign w34[2] = |(datain[303:300] ^ 8);
  assign w34[3] = |(datain[299:296] ^ 14);
  assign w34[4] = |(datain[295:292] ^ 12);
  assign w34[5] = |(datain[291:288] ^ 0);
  assign w34[6] = |(datain[287:284] ^ 11);
  assign w34[7] = |(datain[283:280] ^ 9);
  assign w34[8] = |(datain[279:276] ^ 13);
  assign w34[9] = |(datain[275:272] ^ 8);
  assign w34[10] = |(datain[271:268] ^ 0);
  assign w34[11] = |(datain[267:264] ^ 8);
  assign w34[12] = |(datain[263:260] ^ 11);
  assign w34[13] = |(datain[259:256] ^ 10);
  assign w34[14] = |(datain[255:252] ^ 0);
  assign w34[15] = |(datain[251:248] ^ 0);
  assign w34[16] = |(datain[247:244] ^ 0);
  assign w34[17] = |(datain[243:240] ^ 0);
  assign w34[18] = |(datain[239:236] ^ 14);
  assign w34[19] = |(datain[235:232] ^ 8);
  assign w34[20] = |(datain[231:228] ^ 6);
  assign w34[21] = |(datain[227:224] ^ 10);
  assign w34[22] = |(datain[223:220] ^ 0);
  assign w34[23] = |(datain[219:216] ^ 0);
  assign w34[24] = |(datain[215:212] ^ 5);
  assign w34[25] = |(datain[211:208] ^ 11);
  assign w34[26] = |(datain[207:204] ^ 11);
  assign w34[27] = |(datain[203:200] ^ 4);
  assign w34[28] = |(datain[199:196] ^ 4);
  assign w34[29] = |(datain[195:192] ^ 0);
  assign w34[30] = |(datain[191:188] ^ 12);
  assign w34[31] = |(datain[187:184] ^ 13);
  assign w34[32] = |(datain[183:180] ^ 2);
  assign w34[33] = |(datain[179:176] ^ 1);
  assign w34[34] = |(datain[175:172] ^ 0);
  assign w34[35] = |(datain[171:168] ^ 14);
  assign w34[36] = |(datain[167:164] ^ 1);
  assign w34[37] = |(datain[163:160] ^ 15);
  assign w34[38] = |(datain[159:156] ^ 3);
  assign w34[39] = |(datain[155:152] ^ 3);
  assign w34[40] = |(datain[151:148] ^ 12);
  assign w34[41] = |(datain[147:144] ^ 9);
  assign w34[42] = |(datain[143:140] ^ 3);
  assign w34[43] = |(datain[139:136] ^ 3);
  assign w34[44] = |(datain[135:132] ^ 13);
  assign w34[45] = |(datain[131:128] ^ 2);
  assign w34[46] = |(datain[127:124] ^ 11);
  assign w34[47] = |(datain[123:120] ^ 8);
  assign w34[48] = |(datain[119:116] ^ 0);
  assign w34[49] = |(datain[115:112] ^ 0);
  assign w34[50] = |(datain[111:108] ^ 4);
  assign w34[51] = |(datain[107:104] ^ 2);
  assign w34[52] = |(datain[103:100] ^ 12);
  assign w34[53] = |(datain[99:96] ^ 13);
  assign w34[54] = |(datain[95:92] ^ 2);
  assign w34[55] = |(datain[91:88] ^ 1);
  assign w34[56] = |(datain[87:84] ^ 11);
  assign w34[57] = |(datain[83:80] ^ 4);
  assign w34[58] = |(datain[79:76] ^ 4);
  assign w34[59] = |(datain[75:72] ^ 0);
  assign w34[60] = |(datain[71:68] ^ 11);
  assign w34[61] = |(datain[67:64] ^ 9);
  assign w34[62] = |(datain[63:60] ^ 0);
  assign w34[63] = |(datain[59:56] ^ 4);
  assign w34[64] = |(datain[55:52] ^ 0);
  assign w34[65] = |(datain[51:48] ^ 0);
  assign w34[66] = |(datain[47:44] ^ 11);
  assign w34[67] = |(datain[43:40] ^ 10);
  assign w34[68] = |(datain[39:36] ^ 0);
  assign w34[69] = |(datain[35:32] ^ 2);
  assign w34[70] = |(datain[31:28] ^ 0);
  assign w34[71] = |(datain[27:24] ^ 0);
  assign w34[72] = |(datain[23:20] ^ 12);
  assign w34[73] = |(datain[19:16] ^ 13);
  assign comp[34] = ~(|w34);
  wire [74-1:0] w35;
  assign w35[0] = |(datain[311:308] ^ 4);
  assign w35[1] = |(datain[307:304] ^ 0);
  assign w35[2] = |(datain[303:300] ^ 5);
  assign w35[3] = |(datain[299:296] ^ 9);
  assign w35[4] = |(datain[295:292] ^ 11);
  assign w35[5] = |(datain[291:288] ^ 10);
  assign w35[6] = |(datain[287:284] ^ 3);
  assign w35[7] = |(datain[283:280] ^ 10);
  assign w35[8] = |(datain[279:276] ^ 0);
  assign w35[9] = |(datain[275:272] ^ 4);
  assign w35[10] = |(datain[271:268] ^ 12);
  assign w35[11] = |(datain[267:264] ^ 13);
  assign w35[12] = |(datain[263:260] ^ 2);
  assign w35[13] = |(datain[259:256] ^ 1);
  assign w35[14] = |(datain[255:252] ^ 3);
  assign w35[15] = |(datain[251:248] ^ 2);
  assign w35[16] = |(datain[247:244] ^ 12);
  assign w35[17] = |(datain[243:240] ^ 0);
  assign w35[18] = |(datain[239:236] ^ 14);
  assign w35[19] = |(datain[235:232] ^ 8);
  assign w35[20] = |(datain[231:228] ^ 3);
  assign w35[21] = |(datain[227:224] ^ 1);
  assign w35[22] = |(datain[223:220] ^ 0);
  assign w35[23] = |(datain[219:216] ^ 0);
  assign w35[24] = |(datain[215:212] ^ 11);
  assign w35[25] = |(datain[211:208] ^ 10);
  assign w35[26] = |(datain[207:204] ^ 1);
  assign w35[27] = |(datain[203:200] ^ 11);
  assign w35[28] = |(datain[199:196] ^ 0);
  assign w35[29] = |(datain[195:192] ^ 4);
  assign w35[30] = |(datain[191:188] ^ 12);
  assign w35[31] = |(datain[187:184] ^ 13);
  assign w35[32] = |(datain[183:180] ^ 2);
  assign w35[33] = |(datain[179:176] ^ 1);
  assign w35[34] = |(datain[175:172] ^ 5);
  assign w35[35] = |(datain[171:168] ^ 10);
  assign w35[36] = |(datain[167:164] ^ 5);
  assign w35[37] = |(datain[163:160] ^ 9);
  assign w35[38] = |(datain[159:156] ^ 8);
  assign w35[39] = |(datain[155:152] ^ 0);
  assign w35[40] = |(datain[151:148] ^ 14);
  assign w35[41] = |(datain[147:144] ^ 1);
  assign w35[42] = |(datain[143:140] ^ 14);
  assign w35[43] = |(datain[139:136] ^ 0);
  assign w35[44] = |(datain[135:132] ^ 8);
  assign w35[45] = |(datain[131:128] ^ 0);
  assign w35[46] = |(datain[127:124] ^ 12);
  assign w35[47] = |(datain[123:120] ^ 9);
  assign w35[48] = |(datain[119:116] ^ 0);
  assign w35[49] = |(datain[115:112] ^ 0);
  assign w35[50] = |(datain[111:108] ^ 11);
  assign w35[51] = |(datain[107:104] ^ 8);
  assign w35[52] = |(datain[103:100] ^ 0);
  assign w35[53] = |(datain[99:96] ^ 1);
  assign w35[54] = |(datain[95:92] ^ 5);
  assign w35[55] = |(datain[91:88] ^ 7);
  assign w35[56] = |(datain[87:84] ^ 12);
  assign w35[57] = |(datain[83:80] ^ 13);
  assign w35[58] = |(datain[79:76] ^ 2);
  assign w35[59] = |(datain[75:72] ^ 1);
  assign w35[60] = |(datain[71:68] ^ 1);
  assign w35[61] = |(datain[67:64] ^ 15);
  assign w35[62] = |(datain[63:60] ^ 5);
  assign w35[63] = |(datain[59:56] ^ 10);
  assign w35[64] = |(datain[55:52] ^ 5);
  assign w35[65] = |(datain[51:48] ^ 9);
  assign w35[66] = |(datain[47:44] ^ 14);
  assign w35[67] = |(datain[43:40] ^ 8);
  assign w35[68] = |(datain[39:36] ^ 0);
  assign w35[69] = |(datain[35:32] ^ 15);
  assign w35[70] = |(datain[31:28] ^ 0);
  assign w35[71] = |(datain[27:24] ^ 0);
  assign w35[72] = |(datain[23:20] ^ 11);
  assign w35[73] = |(datain[19:16] ^ 4);
  assign comp[35] = ~(|w35);
  wire [74-1:0] w36;
  assign w36[0] = |(datain[311:308] ^ 3);
  assign w36[1] = |(datain[307:304] ^ 13);
  assign w36[2] = |(datain[303:300] ^ 0);
  assign w36[3] = |(datain[299:296] ^ 7);
  assign w36[4] = |(datain[295:292] ^ 8);
  assign w36[5] = |(datain[291:288] ^ 13);
  assign w36[6] = |(datain[287:284] ^ 11);
  assign w36[7] = |(datain[283:280] ^ 6);
  assign w36[8] = |(datain[279:276] ^ 0);
  assign w36[9] = |(datain[275:272] ^ 8);
  assign w36[10] = |(datain[271:268] ^ 0);
  assign w36[11] = |(datain[267:264] ^ 1);
  assign w36[12] = |(datain[263:260] ^ 14);
  assign w36[13] = |(datain[259:256] ^ 8);
  assign w36[14] = |(datain[255:252] ^ 6);
  assign w36[15] = |(datain[251:248] ^ 8);
  assign w36[16] = |(datain[247:244] ^ 0);
  assign w36[17] = |(datain[243:240] ^ 0);
  assign w36[18] = |(datain[239:236] ^ 8);
  assign w36[19] = |(datain[235:232] ^ 13);
  assign w36[20] = |(datain[231:228] ^ 9);
  assign w36[21] = |(datain[227:224] ^ 6);
  assign w36[22] = |(datain[223:220] ^ 3);
  assign w36[23] = |(datain[219:216] ^ 13);
  assign w36[24] = |(datain[215:212] ^ 0);
  assign w36[25] = |(datain[211:208] ^ 7);
  assign w36[26] = |(datain[207:204] ^ 11);
  assign w36[27] = |(datain[203:200] ^ 4);
  assign w36[28] = |(datain[199:196] ^ 4);
  assign w36[29] = |(datain[195:192] ^ 0);
  assign w36[30] = |(datain[191:188] ^ 12);
  assign w36[31] = |(datain[187:184] ^ 13);
  assign w36[32] = |(datain[183:180] ^ 2);
  assign w36[33] = |(datain[179:176] ^ 1);
  assign w36[34] = |(datain[175:172] ^ 8);
  assign w36[35] = |(datain[171:168] ^ 15);
  assign w36[36] = |(datain[167:164] ^ 8);
  assign w36[37] = |(datain[163:160] ^ 6);
  assign w36[38] = |(datain[159:156] ^ 15);
  assign w36[39] = |(datain[155:152] ^ 15);
  assign w36[40] = |(datain[151:148] ^ 0);
  assign w36[41] = |(datain[147:144] ^ 1);
  assign w36[42] = |(datain[143:140] ^ 11);
  assign w36[43] = |(datain[139:136] ^ 8);
  assign w36[44] = |(datain[135:132] ^ 0);
  assign w36[45] = |(datain[131:128] ^ 0);
  assign w36[46] = |(datain[127:124] ^ 4);
  assign w36[47] = |(datain[123:120] ^ 2);
  assign w36[48] = |(datain[119:116] ^ 14);
  assign w36[49] = |(datain[115:112] ^ 8);
  assign w36[50] = |(datain[111:108] ^ 2);
  assign w36[51] = |(datain[107:104] ^ 11);
  assign w36[52] = |(datain[103:100] ^ 0);
  assign w36[53] = |(datain[99:96] ^ 0);
  assign w36[54] = |(datain[95:92] ^ 8);
  assign w36[55] = |(datain[91:88] ^ 13);
  assign w36[56] = |(datain[87:84] ^ 9);
  assign w36[57] = |(datain[83:80] ^ 6);
  assign w36[58] = |(datain[79:76] ^ 15);
  assign w36[59] = |(datain[75:72] ^ 10);
  assign w36[60] = |(datain[71:68] ^ 0);
  assign w36[61] = |(datain[67:64] ^ 1);
  assign w36[62] = |(datain[63:60] ^ 11);
  assign w36[63] = |(datain[59:56] ^ 9);
  assign w36[64] = |(datain[55:52] ^ 0);
  assign w36[65] = |(datain[51:48] ^ 5);
  assign w36[66] = |(datain[47:44] ^ 0);
  assign w36[67] = |(datain[43:40] ^ 0);
  assign w36[68] = |(datain[39:36] ^ 11);
  assign w36[69] = |(datain[35:32] ^ 4);
  assign w36[70] = |(datain[31:28] ^ 4);
  assign w36[71] = |(datain[27:24] ^ 0);
  assign w36[72] = |(datain[23:20] ^ 12);
  assign w36[73] = |(datain[19:16] ^ 13);
  assign comp[36] = ~(|w36);
  wire [74-1:0] w37;
  assign w37[0] = |(datain[311:308] ^ 11);
  assign w37[1] = |(datain[307:304] ^ 8);
  assign w37[2] = |(datain[303:300] ^ 0);
  assign w37[3] = |(datain[299:296] ^ 0);
  assign w37[4] = |(datain[295:292] ^ 4);
  assign w37[5] = |(datain[291:288] ^ 2);
  assign w37[6] = |(datain[287:284] ^ 14);
  assign w37[7] = |(datain[283:280] ^ 8);
  assign w37[8] = |(datain[279:276] ^ 2);
  assign w37[9] = |(datain[275:272] ^ 11);
  assign w37[10] = |(datain[271:268] ^ 0);
  assign w37[11] = |(datain[267:264] ^ 0);
  assign w37[12] = |(datain[263:260] ^ 8);
  assign w37[13] = |(datain[259:256] ^ 13);
  assign w37[14] = |(datain[255:252] ^ 9);
  assign w37[15] = |(datain[251:248] ^ 6);
  assign w37[16] = |(datain[247:244] ^ 15);
  assign w37[17] = |(datain[243:240] ^ 10);
  assign w37[18] = |(datain[239:236] ^ 0);
  assign w37[19] = |(datain[235:232] ^ 1);
  assign w37[20] = |(datain[231:228] ^ 11);
  assign w37[21] = |(datain[227:224] ^ 9);
  assign w37[22] = |(datain[223:220] ^ 0);
  assign w37[23] = |(datain[219:216] ^ 5);
  assign w37[24] = |(datain[215:212] ^ 0);
  assign w37[25] = |(datain[211:208] ^ 0);
  assign w37[26] = |(datain[207:204] ^ 11);
  assign w37[27] = |(datain[203:200] ^ 4);
  assign w37[28] = |(datain[199:196] ^ 4);
  assign w37[29] = |(datain[195:192] ^ 0);
  assign w37[30] = |(datain[191:188] ^ 12);
  assign w37[31] = |(datain[187:184] ^ 13);
  assign w37[32] = |(datain[183:180] ^ 2);
  assign w37[33] = |(datain[179:176] ^ 1);
  assign w37[34] = |(datain[175:172] ^ 15);
  assign w37[35] = |(datain[171:168] ^ 14);
  assign w37[36] = |(datain[167:164] ^ 8);
  assign w37[37] = |(datain[163:160] ^ 6);
  assign w37[38] = |(datain[159:156] ^ 0);
  assign w37[39] = |(datain[155:152] ^ 1);
  assign w37[40] = |(datain[151:148] ^ 0);
  assign w37[41] = |(datain[147:144] ^ 2);
  assign w37[42] = |(datain[143:140] ^ 5);
  assign w37[43] = |(datain[139:136] ^ 10);
  assign w37[44] = |(datain[135:132] ^ 5);
  assign w37[45] = |(datain[131:128] ^ 9);
  assign w37[46] = |(datain[127:124] ^ 11);
  assign w37[47] = |(datain[123:120] ^ 8);
  assign w37[48] = |(datain[119:116] ^ 0);
  assign w37[49] = |(datain[115:112] ^ 1);
  assign w37[50] = |(datain[111:108] ^ 5);
  assign w37[51] = |(datain[107:104] ^ 7);
  assign w37[52] = |(datain[103:100] ^ 12);
  assign w37[53] = |(datain[99:96] ^ 13);
  assign w37[54] = |(datain[95:92] ^ 2);
  assign w37[55] = |(datain[91:88] ^ 1);
  assign w37[56] = |(datain[87:84] ^ 11);
  assign w37[57] = |(datain[83:80] ^ 4);
  assign w37[58] = |(datain[79:76] ^ 3);
  assign w37[59] = |(datain[75:72] ^ 14);
  assign w37[60] = |(datain[71:68] ^ 12);
  assign w37[61] = |(datain[67:64] ^ 13);
  assign w37[62] = |(datain[63:60] ^ 2);
  assign w37[63] = |(datain[59:56] ^ 1);
  assign w37[64] = |(datain[55:52] ^ 8);
  assign w37[65] = |(datain[51:48] ^ 0);
  assign w37[66] = |(datain[47:44] ^ 11);
  assign w37[67] = |(datain[43:40] ^ 14);
  assign w37[68] = |(datain[39:36] ^ 0);
  assign w37[69] = |(datain[35:32] ^ 1);
  assign w37[70] = |(datain[31:28] ^ 0);
  assign w37[71] = |(datain[27:24] ^ 2);
  assign w37[72] = |(datain[23:20] ^ 0);
  assign w37[73] = |(datain[19:16] ^ 1);
  assign comp[37] = ~(|w37);
  wire [74-1:0] w38;
  assign w38[0] = |(datain[311:308] ^ 15);
  assign w38[1] = |(datain[307:304] ^ 0);
  assign w38[2] = |(datain[303:300] ^ 8);
  assign w38[3] = |(datain[299:296] ^ 11);
  assign w38[4] = |(datain[295:292] ^ 15);
  assign w38[5] = |(datain[291:288] ^ 14);
  assign w38[6] = |(datain[287:284] ^ 11);
  assign w38[7] = |(datain[283:280] ^ 14);
  assign w38[8] = |(datain[279:276] ^ 13);
  assign w38[9] = |(datain[275:272] ^ 2);
  assign w38[10] = |(datain[271:268] ^ 0);
  assign w38[11] = |(datain[267:264] ^ 3);
  assign w38[12] = |(datain[263:260] ^ 11);
  assign w38[13] = |(datain[259:256] ^ 9);
  assign w38[14] = |(datain[255:252] ^ 8);
  assign w38[15] = |(datain[251:248] ^ 6);
  assign w38[16] = |(datain[247:244] ^ 0);
  assign w38[17] = |(datain[243:240] ^ 0);
  assign w38[18] = |(datain[239:236] ^ 15);
  assign w38[19] = |(datain[235:232] ^ 3);
  assign w38[20] = |(datain[231:228] ^ 10);
  assign w38[21] = |(datain[227:224] ^ 4);
  assign w38[22] = |(datain[223:220] ^ 2);
  assign w38[23] = |(datain[219:216] ^ 11);
  assign w38[24] = |(datain[215:212] ^ 13);
  assign w38[25] = |(datain[211:208] ^ 2);
  assign w38[26] = |(datain[207:204] ^ 11);
  assign w38[27] = |(datain[203:200] ^ 9);
  assign w38[28] = |(datain[199:196] ^ 0);
  assign w38[29] = |(datain[195:192] ^ 1);
  assign w38[30] = |(datain[191:188] ^ 0);
  assign w38[31] = |(datain[187:184] ^ 0);
  assign w38[32] = |(datain[183:180] ^ 3);
  assign w38[33] = |(datain[179:176] ^ 2);
  assign w38[34] = |(datain[175:172] ^ 12);
  assign w38[35] = |(datain[171:168] ^ 0);
  assign w38[36] = |(datain[167:164] ^ 11);
  assign w38[37] = |(datain[163:160] ^ 11);
  assign w38[38] = |(datain[159:156] ^ 13);
  assign w38[39] = |(datain[155:152] ^ 8);
  assign w38[40] = |(datain[151:148] ^ 0);
  assign w38[41] = |(datain[147:144] ^ 15);
  assign w38[42] = |(datain[143:140] ^ 12);
  assign w38[43] = |(datain[139:136] ^ 13);
  assign w38[44] = |(datain[135:132] ^ 2);
  assign w38[45] = |(datain[131:128] ^ 6);
  assign w38[46] = |(datain[127:124] ^ 9);
  assign w38[47] = |(datain[123:120] ^ 13);
  assign w38[48] = |(datain[119:116] ^ 7);
  assign w38[49] = |(datain[115:112] ^ 3);
  assign w38[50] = |(datain[111:108] ^ 0);
  assign w38[51] = |(datain[107:104] ^ 3);
  assign w38[52] = |(datain[103:100] ^ 14);
  assign w38[53] = |(datain[99:96] ^ 9);
  assign w38[54] = |(datain[95:92] ^ 6);
  assign w38[55] = |(datain[91:88] ^ 2);
  assign w38[56] = |(datain[87:84] ^ 15);
  assign w38[57] = |(datain[83:80] ^ 14);
  assign w38[58] = |(datain[79:76] ^ 14);
  assign w38[59] = |(datain[75:72] ^ 9);
  assign w38[60] = |(datain[71:68] ^ 6);
  assign w38[61] = |(datain[67:64] ^ 1);
  assign w38[62] = |(datain[63:60] ^ 15);
  assign w38[63] = |(datain[59:56] ^ 14);
  assign w38[64] = |(datain[55:52] ^ 14);
  assign w38[65] = |(datain[51:48] ^ 8);
  assign w38[66] = |(datain[47:44] ^ 0);
  assign w38[67] = |(datain[43:40] ^ 0);
  assign w38[68] = |(datain[39:36] ^ 0);
  assign w38[69] = |(datain[35:32] ^ 0);
  assign w38[70] = |(datain[31:28] ^ 5);
  assign w38[71] = |(datain[27:24] ^ 11);
  assign w38[72] = |(datain[23:20] ^ 8);
  assign w38[73] = |(datain[19:16] ^ 3);
  assign comp[38] = ~(|w38);
  wire [74-1:0] w39;
  assign w39[0] = |(datain[311:308] ^ 2);
  assign w39[1] = |(datain[307:304] ^ 1);
  assign w39[2] = |(datain[303:300] ^ 2);
  assign w39[3] = |(datain[299:296] ^ 6);
  assign w39[4] = |(datain[295:292] ^ 12);
  assign w39[5] = |(datain[291:288] ^ 7);
  assign w39[6] = |(datain[287:284] ^ 4);
  assign w39[7] = |(datain[283:280] ^ 5);
  assign w39[8] = |(datain[279:276] ^ 1);
  assign w39[9] = |(datain[275:272] ^ 5);
  assign w39[10] = |(datain[271:268] ^ 0);
  assign w39[11] = |(datain[267:264] ^ 0);
  assign w39[12] = |(datain[263:260] ^ 0);
  assign w39[13] = |(datain[259:256] ^ 0);
  assign w39[14] = |(datain[255:252] ^ 11);
  assign w39[15] = |(datain[251:248] ^ 4);
  assign w39[16] = |(datain[247:244] ^ 4);
  assign w39[17] = |(datain[243:240] ^ 0);
  assign w39[18] = |(datain[239:236] ^ 11);
  assign w39[19] = |(datain[235:232] ^ 10);
  assign w39[20] = |(datain[231:228] ^ 4);
  assign w39[21] = |(datain[227:224] ^ 9);
  assign w39[22] = |(datain[223:220] ^ 0);
  assign w39[23] = |(datain[219:216] ^ 2);
  assign w39[24] = |(datain[215:212] ^ 11);
  assign w39[25] = |(datain[211:208] ^ 9);
  assign w39[26] = |(datain[207:204] ^ 0);
  assign w39[27] = |(datain[203:200] ^ 5);
  assign w39[28] = |(datain[199:196] ^ 0);
  assign w39[29] = |(datain[195:192] ^ 0);
  assign w39[30] = |(datain[191:188] ^ 12);
  assign w39[31] = |(datain[187:184] ^ 13);
  assign w39[32] = |(datain[183:180] ^ 2);
  assign w39[33] = |(datain[179:176] ^ 1);
  assign w39[34] = |(datain[175:172] ^ 2);
  assign w39[35] = |(datain[171:168] ^ 6);
  assign w39[36] = |(datain[167:164] ^ 8);
  assign w39[37] = |(datain[163:160] ^ 11);
  assign w39[38] = |(datain[159:156] ^ 4);
  assign w39[39] = |(datain[155:152] ^ 13);
  assign w39[40] = |(datain[151:148] ^ 0);
  assign w39[41] = |(datain[147:144] ^ 13);
  assign w39[42] = |(datain[143:140] ^ 2);
  assign w39[43] = |(datain[139:136] ^ 6);
  assign w39[44] = |(datain[135:132] ^ 8);
  assign w39[45] = |(datain[131:128] ^ 11);
  assign w39[46] = |(datain[127:124] ^ 5);
  assign w39[47] = |(datain[123:120] ^ 5);
  assign w39[48] = |(datain[119:116] ^ 0);
  assign w39[49] = |(datain[115:112] ^ 15);
  assign w39[50] = |(datain[111:108] ^ 11);
  assign w39[51] = |(datain[107:104] ^ 8);
  assign w39[52] = |(datain[103:100] ^ 0);
  assign w39[53] = |(datain[99:96] ^ 1);
  assign w39[54] = |(datain[95:92] ^ 5);
  assign w39[55] = |(datain[91:88] ^ 7);
  assign w39[56] = |(datain[87:84] ^ 12);
  assign w39[57] = |(datain[83:80] ^ 13);
  assign w39[58] = |(datain[79:76] ^ 2);
  assign w39[59] = |(datain[75:72] ^ 1);
  assign w39[60] = |(datain[71:68] ^ 11);
  assign w39[61] = |(datain[67:64] ^ 4);
  assign w39[62] = |(datain[63:60] ^ 3);
  assign w39[63] = |(datain[59:56] ^ 14);
  assign w39[64] = |(datain[55:52] ^ 12);
  assign w39[65] = |(datain[51:48] ^ 13);
  assign w39[66] = |(datain[47:44] ^ 2);
  assign w39[67] = |(datain[43:40] ^ 1);
  assign w39[68] = |(datain[39:36] ^ 1);
  assign w39[69] = |(datain[35:32] ^ 15);
  assign w39[70] = |(datain[31:28] ^ 0);
  assign w39[71] = |(datain[27:24] ^ 7);
  assign w39[72] = |(datain[23:20] ^ 5);
  assign w39[73] = |(datain[19:16] ^ 14);
  assign comp[39] = ~(|w39);
  wire [74-1:0] w40;
  assign w40[0] = |(datain[311:308] ^ 0);
  assign w40[1] = |(datain[307:304] ^ 15);
  assign w40[2] = |(datain[303:300] ^ 0);
  assign w40[3] = |(datain[299:296] ^ 0);
  assign w40[4] = |(datain[295:292] ^ 11);
  assign w40[5] = |(datain[291:288] ^ 10);
  assign w40[6] = |(datain[287:284] ^ 13);
  assign w40[7] = |(datain[283:280] ^ 0);
  assign w40[8] = |(datain[279:276] ^ 0);
  assign w40[9] = |(datain[275:272] ^ 9);
  assign w40[10] = |(datain[271:268] ^ 12);
  assign w40[11] = |(datain[267:264] ^ 13);
  assign w40[12] = |(datain[263:260] ^ 2);
  assign w40[13] = |(datain[259:256] ^ 1);
  assign w40[14] = |(datain[255:252] ^ 11);
  assign w40[15] = |(datain[251:248] ^ 8);
  assign w40[16] = |(datain[247:244] ^ 0);
  assign w40[17] = |(datain[243:240] ^ 0);
  assign w40[18] = |(datain[239:236] ^ 4);
  assign w40[19] = |(datain[235:232] ^ 2);
  assign w40[20] = |(datain[231:228] ^ 3);
  assign w40[21] = |(datain[227:224] ^ 3);
  assign w40[22] = |(datain[223:220] ^ 12);
  assign w40[23] = |(datain[219:216] ^ 9);
  assign w40[24] = |(datain[215:212] ^ 9);
  assign w40[25] = |(datain[211:208] ^ 9);
  assign w40[26] = |(datain[207:204] ^ 12);
  assign w40[27] = |(datain[203:200] ^ 13);
  assign w40[28] = |(datain[199:196] ^ 2);
  assign w40[29] = |(datain[195:192] ^ 1);
  assign w40[30] = |(datain[191:188] ^ 11);
  assign w40[31] = |(datain[187:184] ^ 4);
  assign w40[32] = |(datain[183:180] ^ 4);
  assign w40[33] = |(datain[179:176] ^ 0);
  assign w40[34] = |(datain[175:172] ^ 11);
  assign w40[35] = |(datain[171:168] ^ 9);
  assign w40[36] = |(datain[167:164] ^ 2);
  assign w40[37] = |(datain[163:160] ^ 5);
  assign w40[38] = |(datain[159:156] ^ 0);
  assign w40[39] = |(datain[155:152] ^ 0);
  assign w40[40] = |(datain[151:148] ^ 11);
  assign w40[41] = |(datain[147:144] ^ 10);
  assign w40[42] = |(datain[143:140] ^ 14);
  assign w40[43] = |(datain[139:136] ^ 11);
  assign w40[44] = |(datain[135:132] ^ 0);
  assign w40[45] = |(datain[131:128] ^ 8);
  assign w40[46] = |(datain[127:124] ^ 12);
  assign w40[47] = |(datain[123:120] ^ 13);
  assign w40[48] = |(datain[119:116] ^ 2);
  assign w40[49] = |(datain[115:112] ^ 1);
  assign w40[50] = |(datain[111:108] ^ 12);
  assign w40[51] = |(datain[107:104] ^ 3);
  assign w40[52] = |(datain[103:100] ^ 11);
  assign w40[53] = |(datain[99:96] ^ 4);
  assign w40[54] = |(datain[95:92] ^ 4);
  assign w40[55] = |(datain[91:88] ^ 0);
  assign w40[56] = |(datain[87:84] ^ 11);
  assign w40[57] = |(datain[83:80] ^ 9);
  assign w40[58] = |(datain[79:76] ^ 5);
  assign w40[59] = |(datain[75:72] ^ 10);
  assign w40[60] = |(datain[71:68] ^ 0);
  assign w40[61] = |(datain[67:64] ^ 0);
  assign w40[62] = |(datain[63:60] ^ 11);
  assign w40[63] = |(datain[59:56] ^ 10);
  assign w40[64] = |(datain[55:52] ^ 9);
  assign w40[65] = |(datain[51:48] ^ 1);
  assign w40[66] = |(datain[47:44] ^ 0);
  assign w40[67] = |(datain[43:40] ^ 8);
  assign w40[68] = |(datain[39:36] ^ 12);
  assign w40[69] = |(datain[35:32] ^ 13);
  assign w40[70] = |(datain[31:28] ^ 2);
  assign w40[71] = |(datain[27:24] ^ 1);
  assign w40[72] = |(datain[23:20] ^ 5);
  assign w40[73] = |(datain[19:16] ^ 3);
  assign comp[40] = ~(|w40);
  wire [76-1:0] w41;
  assign w41[0] = |(datain[311:308] ^ 12);
  assign w41[1] = |(datain[307:304] ^ 13);
  assign w41[2] = |(datain[303:300] ^ 2);
  assign w41[3] = |(datain[299:296] ^ 1);
  assign w41[4] = |(datain[295:292] ^ 11);
  assign w41[5] = |(datain[291:288] ^ 8);
  assign w41[6] = |(datain[287:284] ^ 0);
  assign w41[7] = |(datain[283:280] ^ 0);
  assign w41[8] = |(datain[279:276] ^ 4);
  assign w41[9] = |(datain[275:272] ^ 2);
  assign w41[10] = |(datain[271:268] ^ 3);
  assign w41[11] = |(datain[267:264] ^ 3);
  assign w41[12] = |(datain[263:260] ^ 12);
  assign w41[13] = |(datain[259:256] ^ 9);
  assign w41[14] = |(datain[255:252] ^ 9);
  assign w41[15] = |(datain[251:248] ^ 9);
  assign w41[16] = |(datain[247:244] ^ 12);
  assign w41[17] = |(datain[243:240] ^ 13);
  assign w41[18] = |(datain[239:236] ^ 2);
  assign w41[19] = |(datain[235:232] ^ 1);
  assign w41[20] = |(datain[231:228] ^ 11);
  assign w41[21] = |(datain[227:224] ^ 10);
  assign w41[22] = |(datain[223:220] ^ 1);
  assign w41[23] = |(datain[219:216] ^ 5);
  assign w41[24] = |(datain[215:212] ^ 0);
  assign w41[25] = |(datain[211:208] ^ 4);
  assign w41[26] = |(datain[207:204] ^ 5);
  assign w41[27] = |(datain[203:200] ^ 9);
  assign w41[28] = |(datain[199:196] ^ 11);
  assign w41[29] = |(datain[195:192] ^ 4);
  assign w41[30] = |(datain[191:188] ^ 4);
  assign w41[31] = |(datain[187:184] ^ 0);
  assign w41[32] = |(datain[183:180] ^ 12);
  assign w41[33] = |(datain[179:176] ^ 13);
  assign w41[34] = |(datain[175:172] ^ 2);
  assign w41[35] = |(datain[171:168] ^ 1);
  assign w41[36] = |(datain[167:164] ^ 11);
  assign w41[37] = |(datain[163:160] ^ 8);
  assign w41[38] = |(datain[159:156] ^ 0);
  assign w41[39] = |(datain[155:152] ^ 1);
  assign w41[40] = |(datain[151:148] ^ 5);
  assign w41[41] = |(datain[147:144] ^ 7);
  assign w41[42] = |(datain[143:140] ^ 5);
  assign w41[43] = |(datain[139:136] ^ 10);
  assign w41[44] = |(datain[135:132] ^ 5);
  assign w41[45] = |(datain[131:128] ^ 9);
  assign w41[46] = |(datain[127:124] ^ 12);
  assign w41[47] = |(datain[123:120] ^ 13);
  assign w41[48] = |(datain[119:116] ^ 2);
  assign w41[49] = |(datain[115:112] ^ 1);
  assign w41[50] = |(datain[111:108] ^ 11);
  assign w41[51] = |(datain[107:104] ^ 4);
  assign w41[52] = |(datain[103:100] ^ 3);
  assign w41[53] = |(datain[99:96] ^ 14);
  assign w41[54] = |(datain[95:92] ^ 12);
  assign w41[55] = |(datain[91:88] ^ 13);
  assign w41[56] = |(datain[87:84] ^ 2);
  assign w41[57] = |(datain[83:80] ^ 1);
  assign w41[58] = |(datain[79:76] ^ 5);
  assign w41[59] = |(datain[75:72] ^ 8);
  assign w41[60] = |(datain[71:68] ^ 5);
  assign w41[61] = |(datain[67:64] ^ 10);
  assign w41[62] = |(datain[63:60] ^ 1);
  assign w41[63] = |(datain[59:56] ^ 15);
  assign w41[64] = |(datain[55:52] ^ 5);
  assign w41[65] = |(datain[51:48] ^ 9);
  assign w41[66] = |(datain[47:44] ^ 12);
  assign w41[67] = |(datain[43:40] ^ 13);
  assign w41[68] = |(datain[39:36] ^ 2);
  assign w41[69] = |(datain[35:32] ^ 1);
  assign w41[70] = |(datain[31:28] ^ 0);
  assign w41[71] = |(datain[27:24] ^ 7);
  assign w41[72] = |(datain[23:20] ^ 1);
  assign w41[73] = |(datain[19:16] ^ 15);
  assign w41[74] = |(datain[15:12] ^ 5);
  assign w41[75] = |(datain[11:8] ^ 15);
  assign comp[41] = ~(|w41);
  wire [76-1:0] w42;
  assign w42[0] = |(datain[311:308] ^ 0);
  assign w42[1] = |(datain[307:304] ^ 4);
  assign w42[2] = |(datain[303:300] ^ 11);
  assign w42[3] = |(datain[299:296] ^ 10);
  assign w42[4] = |(datain[295:292] ^ 0);
  assign w42[5] = |(datain[291:288] ^ 3);
  assign w42[6] = |(datain[287:284] ^ 0);
  assign w42[7] = |(datain[283:280] ^ 1);
  assign w42[8] = |(datain[279:276] ^ 14);
  assign w42[9] = |(datain[275:272] ^ 8);
  assign w42[10] = |(datain[271:268] ^ 9);
  assign w42[11] = |(datain[267:264] ^ 5);
  assign w42[12] = |(datain[263:260] ^ 0);
  assign w42[13] = |(datain[259:256] ^ 1);
  assign w42[14] = |(datain[255:252] ^ 11);
  assign w42[15] = |(datain[251:248] ^ 4);
  assign w42[16] = |(datain[247:244] ^ 4);
  assign w42[17] = |(datain[243:240] ^ 0);
  assign w42[18] = |(datain[239:236] ^ 12);
  assign w42[19] = |(datain[235:232] ^ 13);
  assign w42[20] = |(datain[231:228] ^ 2);
  assign w42[21] = |(datain[227:224] ^ 1);
  assign w42[22] = |(datain[223:220] ^ 0);
  assign w42[23] = |(datain[219:216] ^ 7);
  assign w42[24] = |(datain[215:212] ^ 5);
  assign w42[25] = |(datain[211:208] ^ 15);
  assign w42[26] = |(datain[207:204] ^ 11);
  assign w42[27] = |(datain[203:200] ^ 4);
  assign w42[28] = |(datain[199:196] ^ 4);
  assign w42[29] = |(datain[195:192] ^ 0);
  assign w42[30] = |(datain[191:188] ^ 11);
  assign w42[31] = |(datain[187:184] ^ 9);
  assign w42[32] = |(datain[183:180] ^ 1);
  assign w42[33] = |(datain[179:176] ^ 12);
  assign w42[34] = |(datain[175:172] ^ 0);
  assign w42[35] = |(datain[171:168] ^ 0);
  assign w42[36] = |(datain[167:164] ^ 11);
  assign w42[37] = |(datain[163:160] ^ 10);
  assign w42[38] = |(datain[159:156] ^ 13);
  assign w42[39] = |(datain[155:152] ^ 11);
  assign w42[40] = |(datain[151:148] ^ 0);
  assign w42[41] = |(datain[147:144] ^ 5);
  assign w42[42] = |(datain[143:140] ^ 12);
  assign w42[43] = |(datain[139:136] ^ 13);
  assign w42[44] = |(datain[135:132] ^ 2);
  assign w42[45] = |(datain[131:128] ^ 1);
  assign w42[46] = |(datain[127:124] ^ 14);
  assign w42[47] = |(datain[123:120] ^ 8);
  assign w42[48] = |(datain[119:116] ^ 6);
  assign w42[49] = |(datain[115:112] ^ 12);
  assign w42[50] = |(datain[111:108] ^ 0);
  assign w42[51] = |(datain[107:104] ^ 1);
  assign w42[52] = |(datain[103:100] ^ 11);
  assign w42[53] = |(datain[99:96] ^ 4);
  assign w42[54] = |(datain[95:92] ^ 4);
  assign w42[55] = |(datain[91:88] ^ 0);
  assign w42[56] = |(datain[87:84] ^ 11);
  assign w42[57] = |(datain[83:80] ^ 9);
  assign w42[58] = |(datain[79:76] ^ 1);
  assign w42[59] = |(datain[75:72] ^ 10);
  assign w42[60] = |(datain[71:68] ^ 0);
  assign w42[61] = |(datain[67:64] ^ 0);
  assign w42[62] = |(datain[63:60] ^ 11);
  assign w42[63] = |(datain[59:56] ^ 10);
  assign w42[64] = |(datain[55:52] ^ 3);
  assign w42[65] = |(datain[51:48] ^ 4);
  assign w42[66] = |(datain[47:44] ^ 0);
  assign w42[67] = |(datain[43:40] ^ 11);
  assign w42[68] = |(datain[39:36] ^ 12);
  assign w42[69] = |(datain[35:32] ^ 13);
  assign w42[70] = |(datain[31:28] ^ 2);
  assign w42[71] = |(datain[27:24] ^ 1);
  assign w42[72] = |(datain[23:20] ^ 11);
  assign w42[73] = |(datain[19:16] ^ 8);
  assign w42[74] = |(datain[15:12] ^ 0);
  assign w42[75] = |(datain[11:8] ^ 1);
  assign comp[42] = ~(|w42);
  wire [74-1:0] w43;
  assign w43[0] = |(datain[311:308] ^ 12);
  assign w43[1] = |(datain[307:304] ^ 9);
  assign w43[2] = |(datain[303:300] ^ 8);
  assign w43[3] = |(datain[299:296] ^ 3);
  assign w43[4] = |(datain[295:292] ^ 12);
  assign w43[5] = |(datain[291:288] ^ 2);
  assign w43[6] = |(datain[287:284] ^ 0);
  assign w43[7] = |(datain[283:280] ^ 0);
  assign w43[8] = |(datain[279:276] ^ 11);
  assign w43[9] = |(datain[275:272] ^ 9);
  assign w43[10] = |(datain[271:268] ^ 0);
  assign w43[11] = |(datain[267:264] ^ 4);
  assign w43[12] = |(datain[263:260] ^ 0);
  assign w43[13] = |(datain[259:256] ^ 0);
  assign w43[14] = |(datain[255:252] ^ 8);
  assign w43[15] = |(datain[251:248] ^ 9);
  assign w43[16] = |(datain[247:244] ^ 15);
  assign w43[17] = |(datain[243:240] ^ 15);
  assign w43[18] = |(datain[239:236] ^ 2);
  assign w43[19] = |(datain[235:232] ^ 13);
  assign w43[20] = |(datain[231:228] ^ 0);
  assign w43[21] = |(datain[227:224] ^ 0);
  assign w43[22] = |(datain[223:220] ^ 0);
  assign w43[23] = |(datain[219:216] ^ 0);
  assign w43[24] = |(datain[215:212] ^ 11);
  assign w43[25] = |(datain[211:208] ^ 10);
  assign w43[26] = |(datain[207:204] ^ 3);
  assign w43[27] = |(datain[203:200] ^ 0);
  assign w43[28] = |(datain[199:196] ^ 0);
  assign w43[29] = |(datain[195:192] ^ 1);
  assign w43[30] = |(datain[191:188] ^ 12);
  assign w43[31] = |(datain[187:184] ^ 13);
  assign w43[32] = |(datain[183:180] ^ 2);
  assign w43[33] = |(datain[179:176] ^ 1);
  assign w43[34] = |(datain[175:172] ^ 11);
  assign w43[35] = |(datain[171:168] ^ 8);
  assign w43[36] = |(datain[167:164] ^ 0);
  assign w43[37] = |(datain[163:160] ^ 1);
  assign w43[38] = |(datain[159:156] ^ 5);
  assign w43[39] = |(datain[155:152] ^ 7);
  assign w43[40] = |(datain[151:148] ^ 8);
  assign w43[41] = |(datain[147:144] ^ 11);
  assign w43[42] = |(datain[143:140] ^ 0);
  assign w43[43] = |(datain[139:136] ^ 14);
  assign w43[44] = |(datain[135:132] ^ 4);
  assign w43[45] = |(datain[131:128] ^ 1);
  assign w43[46] = |(datain[127:124] ^ 0);
  assign w43[47] = |(datain[123:120] ^ 1);
  assign w43[48] = |(datain[119:116] ^ 8);
  assign w43[49] = |(datain[115:112] ^ 11);
  assign w43[50] = |(datain[111:108] ^ 1);
  assign w43[51] = |(datain[107:104] ^ 6);
  assign w43[52] = |(datain[103:100] ^ 3);
  assign w43[53] = |(datain[99:96] ^ 15);
  assign w43[54] = |(datain[95:92] ^ 0);
  assign w43[55] = |(datain[91:88] ^ 1);
  assign w43[56] = |(datain[87:84] ^ 8);
  assign w43[57] = |(datain[83:80] ^ 9);
  assign w43[58] = |(datain[79:76] ^ 15);
  assign w43[59] = |(datain[75:72] ^ 15);
  assign w43[60] = |(datain[71:68] ^ 8);
  assign w43[61] = |(datain[67:64] ^ 0);
  assign w43[62] = |(datain[63:60] ^ 12);
  assign w43[63] = |(datain[59:56] ^ 4);
  assign w43[64] = |(datain[55:52] ^ 0);
  assign w43[65] = |(datain[51:48] ^ 0);
  assign w43[66] = |(datain[47:44] ^ 8);
  assign w43[67] = |(datain[43:40] ^ 11);
  assign w43[68] = |(datain[39:36] ^ 1);
  assign w43[69] = |(datain[35:32] ^ 14);
  assign w43[70] = |(datain[31:28] ^ 3);
  assign w43[71] = |(datain[27:24] ^ 6);
  assign w43[72] = |(datain[23:20] ^ 0);
  assign w43[73] = |(datain[19:16] ^ 1);
  assign comp[43] = ~(|w43);
  wire [74-1:0] w44;
  assign w44[0] = |(datain[311:308] ^ 3);
  assign w44[1] = |(datain[307:304] ^ 13);
  assign w44[2] = |(datain[303:300] ^ 11);
  assign w44[3] = |(datain[299:296] ^ 10);
  assign w44[4] = |(datain[295:292] ^ 9);
  assign w44[5] = |(datain[291:288] ^ 14);
  assign w44[6] = |(datain[287:284] ^ 0);
  assign w44[7] = |(datain[283:280] ^ 0);
  assign w44[8] = |(datain[279:276] ^ 12);
  assign w44[9] = |(datain[275:272] ^ 13);
  assign w44[10] = |(datain[271:268] ^ 2);
  assign w44[11] = |(datain[267:264] ^ 1);
  assign w44[12] = |(datain[263:260] ^ 9);
  assign w44[13] = |(datain[259:256] ^ 3);
  assign w44[14] = |(datain[255:252] ^ 11);
  assign w44[15] = |(datain[251:248] ^ 4);
  assign w44[16] = |(datain[247:244] ^ 4);
  assign w44[17] = |(datain[243:240] ^ 0);
  assign w44[18] = |(datain[239:236] ^ 11);
  assign w44[19] = |(datain[235:232] ^ 10);
  assign w44[20] = |(datain[231:228] ^ 0);
  assign w44[21] = |(datain[227:224] ^ 0);
  assign w44[22] = |(datain[223:220] ^ 0);
  assign w44[23] = |(datain[219:216] ^ 1);
  assign w44[24] = |(datain[215:212] ^ 11);
  assign w44[25] = |(datain[211:208] ^ 9);
  assign w44[26] = |(datain[207:204] ^ 13);
  assign w44[27] = |(datain[203:200] ^ 12);
  assign w44[28] = |(datain[199:196] ^ 0);
  assign w44[29] = |(datain[195:192] ^ 0);
  assign w44[30] = |(datain[191:188] ^ 12);
  assign w44[31] = |(datain[187:184] ^ 13);
  assign w44[32] = |(datain[183:180] ^ 2);
  assign w44[33] = |(datain[179:176] ^ 1);
  assign w44[34] = |(datain[175:172] ^ 11);
  assign w44[35] = |(datain[171:168] ^ 4);
  assign w44[36] = |(datain[167:164] ^ 3);
  assign w44[37] = |(datain[163:160] ^ 14);
  assign w44[38] = |(datain[159:156] ^ 12);
  assign w44[39] = |(datain[155:152] ^ 13);
  assign w44[40] = |(datain[151:148] ^ 2);
  assign w44[41] = |(datain[147:144] ^ 1);
  assign w44[42] = |(datain[143:140] ^ 11);
  assign w44[43] = |(datain[139:136] ^ 4);
  assign w44[44] = |(datain[135:132] ^ 4);
  assign w44[45] = |(datain[131:128] ^ 15);
  assign w44[46] = |(datain[127:124] ^ 14);
  assign w44[47] = |(datain[123:120] ^ 9);
  assign w44[48] = |(datain[119:116] ^ 5);
  assign w44[49] = |(datain[115:112] ^ 1);
  assign w44[50] = |(datain[111:108] ^ 15);
  assign w44[51] = |(datain[107:104] ^ 15);
  assign w44[52] = |(datain[103:100] ^ 2);
  assign w44[53] = |(datain[99:96] ^ 10);
  assign w44[54] = |(datain[95:92] ^ 2);
  assign w44[55] = |(datain[91:88] ^ 14);
  assign w44[56] = |(datain[87:84] ^ 6);
  assign w44[57] = |(datain[83:80] ^ 5);
  assign w44[58] = |(datain[79:76] ^ 7);
  assign w44[59] = |(datain[75:72] ^ 8);
  assign w44[60] = |(datain[71:68] ^ 6);
  assign w44[61] = |(datain[67:64] ^ 5);
  assign w44[62] = |(datain[63:60] ^ 0);
  assign w44[63] = |(datain[59:56] ^ 0);
  assign w44[64] = |(datain[55:52] ^ 5);
  assign w44[65] = |(datain[51:48] ^ 11);
  assign w44[66] = |(datain[47:44] ^ 4);
  assign w44[67] = |(datain[43:40] ^ 12);
  assign w44[68] = |(datain[39:36] ^ 6);
  assign w44[69] = |(datain[35:32] ^ 9);
  assign w44[70] = |(datain[31:28] ^ 7);
  assign w44[71] = |(datain[27:24] ^ 6);
  assign w44[72] = |(datain[23:20] ^ 6);
  assign w44[73] = |(datain[19:16] ^ 5);
  assign comp[44] = ~(|w44);
  wire [76-1:0] w45;
  assign w45[0] = |(datain[311:308] ^ 12);
  assign w45[1] = |(datain[307:304] ^ 9);
  assign w45[2] = |(datain[303:300] ^ 11);
  assign w45[3] = |(datain[299:296] ^ 8);
  assign w45[4] = |(datain[295:292] ^ 0);
  assign w45[5] = |(datain[291:288] ^ 0);
  assign w45[6] = |(datain[287:284] ^ 4);
  assign w45[7] = |(datain[283:280] ^ 2);
  assign w45[8] = |(datain[279:276] ^ 3);
  assign w45[9] = |(datain[275:272] ^ 3);
  assign w45[10] = |(datain[271:268] ^ 13);
  assign w45[11] = |(datain[267:264] ^ 2);
  assign w45[12] = |(datain[263:260] ^ 12);
  assign w45[13] = |(datain[259:256] ^ 13);
  assign w45[14] = |(datain[255:252] ^ 2);
  assign w45[15] = |(datain[251:248] ^ 1);
  assign w45[16] = |(datain[247:244] ^ 11);
  assign w45[17] = |(datain[243:240] ^ 4);
  assign w45[18] = |(datain[239:236] ^ 4);
  assign w45[19] = |(datain[235:232] ^ 0);
  assign w45[20] = |(datain[231:228] ^ 11);
  assign w45[21] = |(datain[227:224] ^ 9);
  assign w45[22] = |(datain[223:220] ^ 0);
  assign w45[23] = |(datain[219:216] ^ 3);
  assign w45[24] = |(datain[215:212] ^ 0);
  assign w45[25] = |(datain[211:208] ^ 0);
  assign w45[26] = |(datain[207:204] ^ 11);
  assign w45[27] = |(datain[203:200] ^ 10);
  assign w45[28] = |(datain[199:196] ^ 7);
  assign w45[29] = |(datain[195:192] ^ 7);
  assign w45[30] = |(datain[191:188] ^ 0);
  assign w45[31] = |(datain[187:184] ^ 3);
  assign w45[32] = |(datain[183:180] ^ 12);
  assign w45[33] = |(datain[179:176] ^ 13);
  assign w45[34] = |(datain[175:172] ^ 2);
  assign w45[35] = |(datain[171:168] ^ 1);
  assign w45[36] = |(datain[167:164] ^ 11);
  assign w45[37] = |(datain[163:160] ^ 8);
  assign w45[38] = |(datain[159:156] ^ 0);
  assign w45[39] = |(datain[155:152] ^ 1);
  assign w45[40] = |(datain[151:148] ^ 5);
  assign w45[41] = |(datain[147:144] ^ 7);
  assign w45[42] = |(datain[143:140] ^ 5);
  assign w45[43] = |(datain[139:136] ^ 10);
  assign w45[44] = |(datain[135:132] ^ 5);
  assign w45[45] = |(datain[131:128] ^ 9);
  assign w45[46] = |(datain[127:124] ^ 12);
  assign w45[47] = |(datain[123:120] ^ 13);
  assign w45[48] = |(datain[119:116] ^ 2);
  assign w45[49] = |(datain[115:112] ^ 1);
  assign w45[50] = |(datain[111:108] ^ 11);
  assign w45[51] = |(datain[107:104] ^ 4);
  assign w45[52] = |(datain[103:100] ^ 3);
  assign w45[53] = |(datain[99:96] ^ 14);
  assign w45[54] = |(datain[95:92] ^ 12);
  assign w45[55] = |(datain[91:88] ^ 13);
  assign w45[56] = |(datain[87:84] ^ 2);
  assign w45[57] = |(datain[83:80] ^ 1);
  assign w45[58] = |(datain[79:76] ^ 5);
  assign w45[59] = |(datain[75:72] ^ 8);
  assign w45[60] = |(datain[71:68] ^ 5);
  assign w45[61] = |(datain[67:64] ^ 10);
  assign w45[62] = |(datain[63:60] ^ 1);
  assign w45[63] = |(datain[59:56] ^ 15);
  assign w45[64] = |(datain[55:52] ^ 5);
  assign w45[65] = |(datain[51:48] ^ 9);
  assign w45[66] = |(datain[47:44] ^ 12);
  assign w45[67] = |(datain[43:40] ^ 13);
  assign w45[68] = |(datain[39:36] ^ 2);
  assign w45[69] = |(datain[35:32] ^ 1);
  assign w45[70] = |(datain[31:28] ^ 5);
  assign w45[71] = |(datain[27:24] ^ 10);
  assign w45[72] = |(datain[23:20] ^ 1);
  assign w45[73] = |(datain[19:16] ^ 15);
  assign w45[74] = |(datain[15:12] ^ 11);
  assign w45[75] = |(datain[11:8] ^ 8);
  assign comp[45] = ~(|w45);
  wire [76-1:0] w46;
  assign w46[0] = |(datain[311:308] ^ 12);
  assign w46[1] = |(datain[307:304] ^ 13);
  assign w46[2] = |(datain[303:300] ^ 2);
  assign w46[3] = |(datain[299:296] ^ 1);
  assign w46[4] = |(datain[295:292] ^ 8);
  assign w46[5] = |(datain[291:288] ^ 0);
  assign w46[6] = |(datain[287:284] ^ 15);
  assign w46[7] = |(datain[283:280] ^ 10);
  assign w46[8] = |(datain[279:276] ^ 0);
  assign w46[9] = |(datain[275:272] ^ 0);
  assign w46[10] = |(datain[271:268] ^ 7);
  assign w46[11] = |(datain[267:264] ^ 5);
  assign w46[12] = |(datain[263:260] ^ 1);
  assign w46[13] = |(datain[259:256] ^ 5);
  assign w46[14] = |(datain[255:252] ^ 11);
  assign w46[15] = |(datain[251:248] ^ 8);
  assign w46[16] = |(datain[247:244] ^ 0);
  assign w46[17] = |(datain[243:240] ^ 2);
  assign w46[18] = |(datain[239:236] ^ 4);
  assign w46[19] = |(datain[235:232] ^ 2);
  assign w46[20] = |(datain[231:228] ^ 3);
  assign w46[21] = |(datain[227:224] ^ 3);
  assign w46[22] = |(datain[223:220] ^ 12);
  assign w46[23] = |(datain[219:216] ^ 9);
  assign w46[24] = |(datain[215:212] ^ 3);
  assign w46[25] = |(datain[211:208] ^ 3);
  assign w46[26] = |(datain[207:204] ^ 13);
  assign w46[27] = |(datain[203:200] ^ 2);
  assign w46[28] = |(datain[199:196] ^ 12);
  assign w46[29] = |(datain[195:192] ^ 13);
  assign w46[30] = |(datain[191:188] ^ 2);
  assign w46[31] = |(datain[187:184] ^ 1);
  assign w46[32] = |(datain[183:180] ^ 0);
  assign w46[33] = |(datain[179:176] ^ 14);
  assign w46[34] = |(datain[175:172] ^ 1);
  assign w46[35] = |(datain[171:168] ^ 15);
  assign w46[36] = |(datain[167:164] ^ 11);
  assign w46[37] = |(datain[163:160] ^ 4);
  assign w46[38] = |(datain[159:156] ^ 4);
  assign w46[39] = |(datain[155:152] ^ 0);
  assign w46[40] = |(datain[151:148] ^ 11);
  assign w46[41] = |(datain[147:144] ^ 10);
  assign w46[42] = |(datain[143:140] ^ 10);
  assign w46[43] = |(datain[139:136] ^ 5);
  assign w46[44] = |(datain[135:132] ^ 0);
  assign w46[45] = |(datain[131:128] ^ 2);
  assign w46[46] = |(datain[127:124] ^ 11);
  assign w46[47] = |(datain[123:120] ^ 9);
  assign w46[48] = |(datain[119:116] ^ 1);
  assign w46[49] = |(datain[115:112] ^ 13);
  assign w46[50] = |(datain[111:108] ^ 0);
  assign w46[51] = |(datain[107:104] ^ 0);
  assign w46[52] = |(datain[103:100] ^ 12);
  assign w46[53] = |(datain[99:96] ^ 13);
  assign w46[54] = |(datain[95:92] ^ 2);
  assign w46[55] = |(datain[91:88] ^ 1);
  assign w46[56] = |(datain[87:84] ^ 0);
  assign w46[57] = |(datain[83:80] ^ 14);
  assign w46[58] = |(datain[79:76] ^ 1);
  assign w46[59] = |(datain[75:72] ^ 15);
  assign w46[60] = |(datain[71:68] ^ 11);
  assign w46[61] = |(datain[67:64] ^ 8);
  assign w46[62] = |(datain[63:60] ^ 0);
  assign w46[63] = |(datain[59:56] ^ 1);
  assign w46[64] = |(datain[55:52] ^ 5);
  assign w46[65] = |(datain[51:48] ^ 7);
  assign w46[66] = |(datain[47:44] ^ 8);
  assign w46[67] = |(datain[43:40] ^ 11);
  assign w46[68] = |(datain[39:36] ^ 0);
  assign w46[69] = |(datain[35:32] ^ 14);
  assign w46[70] = |(datain[31:28] ^ 10);
  assign w46[71] = |(datain[27:24] ^ 1);
  assign w46[72] = |(datain[23:20] ^ 0);
  assign w46[73] = |(datain[19:16] ^ 2);
  assign w46[74] = |(datain[15:12] ^ 8);
  assign w46[75] = |(datain[11:8] ^ 11);
  assign comp[46] = ~(|w46);
  wire [76-1:0] w47;
  assign w47[0] = |(datain[311:308] ^ 12);
  assign w47[1] = |(datain[307:304] ^ 13);
  assign w47[2] = |(datain[303:300] ^ 2);
  assign w47[3] = |(datain[299:296] ^ 1);
  assign w47[4] = |(datain[295:292] ^ 15);
  assign w47[5] = |(datain[291:288] ^ 14);
  assign w47[6] = |(datain[287:284] ^ 12);
  assign w47[7] = |(datain[283:280] ^ 0);
  assign w47[8] = |(datain[279:276] ^ 13);
  assign w47[9] = |(datain[275:272] ^ 0);
  assign w47[10] = |(datain[271:268] ^ 14);
  assign w47[11] = |(datain[267:264] ^ 0);
  assign w47[12] = |(datain[263:260] ^ 3);
  assign w47[13] = |(datain[259:256] ^ 10);
  assign w47[14] = |(datain[255:252] ^ 13);
  assign w47[15] = |(datain[251:248] ^ 0);
  assign w47[16] = |(datain[247:244] ^ 7);
  assign w47[17] = |(datain[243:240] ^ 5);
  assign w47[18] = |(datain[239:236] ^ 3);
  assign w47[19] = |(datain[235:232] ^ 3);
  assign w47[20] = |(datain[231:228] ^ 11);
  assign w47[21] = |(datain[227:224] ^ 4);
  assign w47[22] = |(datain[223:220] ^ 1);
  assign w47[23] = |(datain[219:216] ^ 3);
  assign w47[24] = |(datain[215:212] ^ 12);
  assign w47[25] = |(datain[211:208] ^ 13);
  assign w47[26] = |(datain[207:204] ^ 2);
  assign w47[27] = |(datain[203:200] ^ 15);
  assign w47[28] = |(datain[199:196] ^ 1);
  assign w47[29] = |(datain[195:192] ^ 14);
  assign w47[30] = |(datain[191:188] ^ 5);
  assign w47[31] = |(datain[187:184] ^ 2);
  assign w47[32] = |(datain[183:180] ^ 11);
  assign w47[33] = |(datain[179:176] ^ 4);
  assign w47[34] = |(datain[175:172] ^ 1);
  assign w47[35] = |(datain[171:168] ^ 3);
  assign w47[36] = |(datain[167:164] ^ 12);
  assign w47[37] = |(datain[163:160] ^ 13);
  assign w47[38] = |(datain[159:156] ^ 2);
  assign w47[39] = |(datain[155:152] ^ 15);
  assign w47[40] = |(datain[151:148] ^ 5);
  assign w47[41] = |(datain[147:144] ^ 10);
  assign w47[42] = |(datain[143:140] ^ 1);
  assign w47[43] = |(datain[139:136] ^ 15);
  assign w47[44] = |(datain[135:132] ^ 11);
  assign w47[45] = |(datain[131:128] ^ 8);
  assign w47[46] = |(datain[127:124] ^ 1);
  assign w47[47] = |(datain[123:120] ^ 3);
  assign w47[48] = |(datain[119:116] ^ 2);
  assign w47[49] = |(datain[115:112] ^ 5);
  assign w47[50] = |(datain[111:108] ^ 12);
  assign w47[51] = |(datain[107:104] ^ 13);
  assign w47[52] = |(datain[103:100] ^ 2);
  assign w47[53] = |(datain[99:96] ^ 1);
  assign w47[54] = |(datain[95:92] ^ 11);
  assign w47[55] = |(datain[91:88] ^ 9);
  assign w47[56] = |(datain[87:84] ^ 0);
  assign w47[57] = |(datain[83:80] ^ 1);
  assign w47[58] = |(datain[79:76] ^ 0);
  assign w47[59] = |(datain[75:72] ^ 0);
  assign w47[60] = |(datain[71:68] ^ 11);
  assign w47[61] = |(datain[67:64] ^ 10);
  assign w47[62] = |(datain[63:60] ^ 8);
  assign w47[63] = |(datain[59:56] ^ 0);
  assign w47[64] = |(datain[55:52] ^ 0);
  assign w47[65] = |(datain[51:48] ^ 5);
  assign w47[66] = |(datain[47:44] ^ 11);
  assign w47[67] = |(datain[43:40] ^ 8);
  assign w47[68] = |(datain[39:36] ^ 0);
  assign w47[69] = |(datain[35:32] ^ 8);
  assign w47[70] = |(datain[31:28] ^ 0);
  assign w47[71] = |(datain[27:24] ^ 3);
  assign w47[72] = |(datain[23:20] ^ 12);
  assign w47[73] = |(datain[19:16] ^ 13);
  assign w47[74] = |(datain[15:12] ^ 1);
  assign w47[75] = |(datain[11:8] ^ 3);
  assign comp[47] = ~(|w47);
  wire [76-1:0] w48;
  assign w48[0] = |(datain[311:308] ^ 2);
  assign w48[1] = |(datain[307:304] ^ 13);
  assign w48[2] = |(datain[303:300] ^ 0);
  assign w48[3] = |(datain[299:296] ^ 4);
  assign w48[4] = |(datain[295:292] ^ 0);
  assign w48[5] = |(datain[291:288] ^ 0);
  assign w48[6] = |(datain[287:284] ^ 2);
  assign w48[7] = |(datain[283:280] ^ 14);
  assign w48[8] = |(datain[279:276] ^ 8);
  assign w48[9] = |(datain[275:272] ^ 9);
  assign w48[10] = |(datain[271:268] ^ 8);
  assign w48[11] = |(datain[267:264] ^ 6);
  assign w48[12] = |(datain[263:260] ^ 1);
  assign w48[13] = |(datain[259:256] ^ 7);
  assign w48[14] = |(datain[255:252] ^ 0);
  assign w48[15] = |(datain[251:248] ^ 1);
  assign w48[16] = |(datain[247:244] ^ 11);
  assign w48[17] = |(datain[243:240] ^ 4);
  assign w48[18] = |(datain[239:236] ^ 4);
  assign w48[19] = |(datain[235:232] ^ 0);
  assign w48[20] = |(datain[231:228] ^ 8);
  assign w48[21] = |(datain[227:224] ^ 11);
  assign w48[22] = |(datain[223:220] ^ 13);
  assign w48[23] = |(datain[219:216] ^ 5);
  assign w48[24] = |(datain[215:212] ^ 11);
  assign w48[25] = |(datain[211:208] ^ 9);
  assign w48[26] = |(datain[207:204] ^ 5);
  assign w48[27] = |(datain[203:200] ^ 7);
  assign w48[28] = |(datain[199:196] ^ 0);
  assign w48[29] = |(datain[195:192] ^ 1);
  assign w48[30] = |(datain[191:188] ^ 9);
  assign w48[31] = |(datain[187:184] ^ 0);
  assign w48[32] = |(datain[183:180] ^ 12);
  assign w48[33] = |(datain[179:176] ^ 13);
  assign w48[34] = |(datain[175:172] ^ 2);
  assign w48[35] = |(datain[171:168] ^ 1);
  assign w48[36] = |(datain[167:164] ^ 11);
  assign w48[37] = |(datain[163:160] ^ 8);
  assign w48[38] = |(datain[159:156] ^ 0);
  assign w48[39] = |(datain[155:152] ^ 0);
  assign w48[40] = |(datain[151:148] ^ 4);
  assign w48[41] = |(datain[147:144] ^ 2);
  assign w48[42] = |(datain[143:140] ^ 3);
  assign w48[43] = |(datain[139:136] ^ 3);
  assign w48[44] = |(datain[135:132] ^ 12);
  assign w48[45] = |(datain[131:128] ^ 9);
  assign w48[46] = |(datain[127:124] ^ 3);
  assign w48[47] = |(datain[123:120] ^ 3);
  assign w48[48] = |(datain[119:116] ^ 13);
  assign w48[49] = |(datain[115:112] ^ 2);
  assign w48[50] = |(datain[111:108] ^ 12);
  assign w48[51] = |(datain[107:104] ^ 13);
  assign w48[52] = |(datain[103:100] ^ 2);
  assign w48[53] = |(datain[99:96] ^ 1);
  assign w48[54] = |(datain[95:92] ^ 11);
  assign w48[55] = |(datain[91:88] ^ 4);
  assign w48[56] = |(datain[87:84] ^ 4);
  assign w48[57] = |(datain[83:80] ^ 0);
  assign w48[58] = |(datain[79:76] ^ 8);
  assign w48[59] = |(datain[75:72] ^ 11);
  assign w48[60] = |(datain[71:68] ^ 13);
  assign w48[61] = |(datain[67:64] ^ 5);
  assign w48[62] = |(datain[63:60] ^ 8);
  assign w48[63] = |(datain[59:56] ^ 1);
  assign w48[64] = |(datain[55:52] ^ 12);
  assign w48[65] = |(datain[51:48] ^ 2);
  assign w48[66] = |(datain[47:44] ^ 1);
  assign w48[67] = |(datain[43:40] ^ 5);
  assign w48[68] = |(datain[39:36] ^ 0);
  assign w48[69] = |(datain[35:32] ^ 1);
  assign w48[70] = |(datain[31:28] ^ 11);
  assign w48[71] = |(datain[27:24] ^ 9);
  assign w48[72] = |(datain[23:20] ^ 0);
  assign w48[73] = |(datain[19:16] ^ 4);
  assign w48[74] = |(datain[15:12] ^ 0);
  assign w48[75] = |(datain[11:8] ^ 0);
  assign comp[48] = ~(|w48);
  wire [76-1:0] w49;
  assign w49[0] = |(datain[311:308] ^ 14);
  assign w49[1] = |(datain[307:304] ^ 8);
  assign w49[2] = |(datain[303:300] ^ 1);
  assign w49[3] = |(datain[299:296] ^ 2);
  assign w49[4] = |(datain[295:292] ^ 0);
  assign w49[5] = |(datain[291:288] ^ 0);
  assign w49[6] = |(datain[287:284] ^ 4);
  assign w49[7] = |(datain[283:280] ^ 8);
  assign w49[8] = |(datain[279:276] ^ 4);
  assign w49[9] = |(datain[275:272] ^ 8);
  assign w49[10] = |(datain[271:268] ^ 4);
  assign w49[11] = |(datain[267:264] ^ 8);
  assign w49[12] = |(datain[263:260] ^ 10);
  assign w49[13] = |(datain[259:256] ^ 3);
  assign w49[14] = |(datain[255:252] ^ 6);
  assign w49[15] = |(datain[251:248] ^ 7);
  assign w49[16] = |(datain[247:244] ^ 0);
  assign w49[17] = |(datain[243:240] ^ 0);
  assign w49[18] = |(datain[239:236] ^ 5);
  assign w49[19] = |(datain[235:232] ^ 3);
  assign w49[20] = |(datain[231:228] ^ 14);
  assign w49[21] = |(datain[227:224] ^ 8);
  assign w49[22] = |(datain[223:220] ^ 8);
  assign w49[23] = |(datain[219:216] ^ 0);
  assign w49[24] = |(datain[215:212] ^ 0);
  assign w49[25] = |(datain[211:208] ^ 0);
  assign w49[26] = |(datain[207:204] ^ 5);
  assign w49[27] = |(datain[203:200] ^ 11);
  assign w49[28] = |(datain[199:196] ^ 11);
  assign w49[29] = |(datain[195:192] ^ 4);
  assign w49[30] = |(datain[191:188] ^ 4);
  assign w49[31] = |(datain[187:184] ^ 0);
  assign w49[32] = |(datain[183:180] ^ 12);
  assign w49[33] = |(datain[179:176] ^ 13);
  assign w49[34] = |(datain[175:172] ^ 2);
  assign w49[35] = |(datain[171:168] ^ 1);
  assign w49[36] = |(datain[167:164] ^ 11);
  assign w49[37] = |(datain[163:160] ^ 8);
  assign w49[38] = |(datain[159:156] ^ 0);
  assign w49[39] = |(datain[155:152] ^ 0);
  assign w49[40] = |(datain[151:148] ^ 4);
  assign w49[41] = |(datain[147:144] ^ 2);
  assign w49[42] = |(datain[143:140] ^ 9);
  assign w49[43] = |(datain[139:136] ^ 9);
  assign w49[44] = |(datain[135:132] ^ 3);
  assign w49[45] = |(datain[131:128] ^ 3);
  assign w49[46] = |(datain[127:124] ^ 12);
  assign w49[47] = |(datain[123:120] ^ 9);
  assign w49[48] = |(datain[119:116] ^ 12);
  assign w49[49] = |(datain[115:112] ^ 13);
  assign w49[50] = |(datain[111:108] ^ 2);
  assign w49[51] = |(datain[107:104] ^ 1);
  assign w49[52] = |(datain[103:100] ^ 12);
  assign w49[53] = |(datain[99:96] ^ 3);
  assign w49[54] = |(datain[95:92] ^ 12);
  assign w49[55] = |(datain[91:88] ^ 3);
  assign w49[56] = |(datain[87:84] ^ 12);
  assign w49[57] = |(datain[83:80] ^ 3);
  assign w49[58] = |(datain[79:76] ^ 3);
  assign w49[59] = |(datain[75:72] ^ 13);
  assign w49[60] = |(datain[71:68] ^ 0);
  assign w49[61] = |(datain[67:64] ^ 0);
  assign w49[62] = |(datain[63:60] ^ 4);
  assign w49[63] = |(datain[59:56] ^ 11);
  assign w49[64] = |(datain[55:52] ^ 5);
  assign w49[65] = |(datain[51:48] ^ 0);
  assign w49[66] = |(datain[47:44] ^ 5);
  assign w49[67] = |(datain[43:40] ^ 3);
  assign w49[68] = |(datain[39:36] ^ 7);
  assign w49[69] = |(datain[35:32] ^ 5);
  assign w49[70] = |(datain[31:28] ^ 6);
  assign w49[71] = |(datain[27:24] ^ 5);
  assign w49[72] = |(datain[23:20] ^ 11);
  assign w49[73] = |(datain[19:16] ^ 4);
  assign w49[74] = |(datain[15:12] ^ 4);
  assign w49[75] = |(datain[11:8] ^ 3);
  assign comp[49] = ~(|w49);
  wire [76-1:0] w50;
  assign w50[0] = |(datain[311:308] ^ 0);
  assign w50[1] = |(datain[307:304] ^ 3);
  assign w50[2] = |(datain[303:300] ^ 11);
  assign w50[3] = |(datain[299:296] ^ 15);
  assign w50[4] = |(datain[295:292] ^ 11);
  assign w50[5] = |(datain[291:288] ^ 2);
  assign w50[6] = |(datain[287:284] ^ 0);
  assign w50[7] = |(datain[283:280] ^ 3);
  assign w50[8] = |(datain[279:276] ^ 5);
  assign w50[9] = |(datain[275:272] ^ 7);
  assign w50[10] = |(datain[271:268] ^ 3);
  assign w50[11] = |(datain[267:264] ^ 3);
  assign w50[12] = |(datain[263:260] ^ 15);
  assign w50[13] = |(datain[259:256] ^ 6);
  assign w50[14] = |(datain[255:252] ^ 8);
  assign w50[15] = |(datain[251:248] ^ 1);
  assign w50[16] = |(datain[247:244] ^ 12);
  assign w50[17] = |(datain[243:240] ^ 5);
  assign w50[18] = |(datain[239:236] ^ 0);
  assign w50[19] = |(datain[235:232] ^ 0);
  assign w50[20] = |(datain[231:228] ^ 0);
  assign w50[21] = |(datain[227:224] ^ 1);
  assign w50[22] = |(datain[223:220] ^ 14);
  assign w50[23] = |(datain[219:216] ^ 8);
  assign w50[24] = |(datain[215:212] ^ 8);
  assign w50[25] = |(datain[211:208] ^ 7);
  assign w50[26] = |(datain[207:204] ^ 0);
  assign w50[27] = |(datain[203:200] ^ 1);
  assign w50[28] = |(datain[199:196] ^ 11);
  assign w50[29] = |(datain[195:192] ^ 4);
  assign w50[30] = |(datain[191:188] ^ 4);
  assign w50[31] = |(datain[187:184] ^ 0);
  assign w50[32] = |(datain[183:180] ^ 11);
  assign w50[33] = |(datain[179:176] ^ 9);
  assign w50[34] = |(datain[175:172] ^ 12);
  assign w50[35] = |(datain[171:168] ^ 1);
  assign w50[36] = |(datain[167:164] ^ 0);
  assign w50[37] = |(datain[163:160] ^ 4);
  assign w50[38] = |(datain[159:156] ^ 5);
  assign w50[39] = |(datain[155:152] ^ 10);
  assign w50[40] = |(datain[151:148] ^ 12);
  assign w50[41] = |(datain[147:144] ^ 13);
  assign w50[42] = |(datain[143:140] ^ 2);
  assign w50[43] = |(datain[139:136] ^ 1);
  assign w50[44] = |(datain[135:132] ^ 11);
  assign w50[45] = |(datain[131:128] ^ 8);
  assign w50[46] = |(datain[127:124] ^ 0);
  assign w50[47] = |(datain[123:120] ^ 0);
  assign w50[48] = |(datain[119:116] ^ 4);
  assign w50[49] = |(datain[115:112] ^ 2);
  assign w50[50] = |(datain[111:108] ^ 14);
  assign w50[51] = |(datain[107:104] ^ 8);
  assign w50[52] = |(datain[103:100] ^ 4);
  assign w50[53] = |(datain[99:96] ^ 0);
  assign w50[54] = |(datain[95:92] ^ 0);
  assign w50[55] = |(datain[91:88] ^ 0);
  assign w50[56] = |(datain[87:84] ^ 11);
  assign w50[57] = |(datain[83:80] ^ 4);
  assign w50[58] = |(datain[79:76] ^ 4);
  assign w50[59] = |(datain[75:72] ^ 0);
  assign w50[60] = |(datain[71:68] ^ 11);
  assign w50[61] = |(datain[67:64] ^ 9);
  assign w50[62] = |(datain[63:60] ^ 0);
  assign w50[63] = |(datain[59:56] ^ 4);
  assign w50[64] = |(datain[55:52] ^ 0);
  assign w50[65] = |(datain[51:48] ^ 0);
  assign w50[66] = |(datain[47:44] ^ 11);
  assign w50[67] = |(datain[43:40] ^ 10);
  assign w50[68] = |(datain[39:36] ^ 2);
  assign w50[69] = |(datain[35:32] ^ 0);
  assign w50[70] = |(datain[31:28] ^ 0);
  assign w50[71] = |(datain[27:24] ^ 3);
  assign w50[72] = |(datain[23:20] ^ 12);
  assign w50[73] = |(datain[19:16] ^ 13);
  assign w50[74] = |(datain[15:12] ^ 2);
  assign w50[75] = |(datain[11:8] ^ 1);
  assign comp[50] = ~(|w50);
  wire [74-1:0] w51;
  assign w51[0] = |(datain[311:308] ^ 14);
  assign w51[1] = |(datain[307:304] ^ 8);
  assign w51[2] = |(datain[303:300] ^ 8);
  assign w51[3] = |(datain[299:296] ^ 12);
  assign w51[4] = |(datain[295:292] ^ 0);
  assign w51[5] = |(datain[291:288] ^ 0);
  assign w51[6] = |(datain[287:284] ^ 11);
  assign w51[7] = |(datain[283:280] ^ 0);
  assign w51[8] = |(datain[279:276] ^ 0);
  assign w51[9] = |(datain[275:272] ^ 2);
  assign w51[10] = |(datain[271:268] ^ 14);
  assign w51[11] = |(datain[267:264] ^ 8);
  assign w51[12] = |(datain[263:260] ^ 7);
  assign w51[13] = |(datain[259:256] ^ 13);
  assign w51[14] = |(datain[255:252] ^ 0);
  assign w51[15] = |(datain[251:248] ^ 0);
  assign w51[16] = |(datain[247:244] ^ 11);
  assign w51[17] = |(datain[243:240] ^ 4);
  assign w51[18] = |(datain[239:236] ^ 4);
  assign w51[19] = |(datain[235:232] ^ 0);
  assign w51[20] = |(datain[231:228] ^ 8);
  assign w51[21] = |(datain[227:224] ^ 13);
  assign w51[22] = |(datain[223:220] ^ 9);
  assign w51[23] = |(datain[219:216] ^ 6);
  assign w51[24] = |(datain[215:212] ^ 4);
  assign w51[25] = |(datain[211:208] ^ 7);
  assign w51[26] = |(datain[207:204] ^ 0);
  assign w51[27] = |(datain[203:200] ^ 3);
  assign w51[28] = |(datain[199:196] ^ 5);
  assign w51[29] = |(datain[195:192] ^ 9);
  assign w51[30] = |(datain[191:188] ^ 12);
  assign w51[31] = |(datain[187:184] ^ 13);
  assign w51[32] = |(datain[183:180] ^ 2);
  assign w51[33] = |(datain[179:176] ^ 1);
  assign w51[34] = |(datain[175:172] ^ 11);
  assign w51[35] = |(datain[171:168] ^ 8);
  assign w51[36] = |(datain[167:164] ^ 0);
  assign w51[37] = |(datain[163:160] ^ 2);
  assign w51[38] = |(datain[159:156] ^ 4);
  assign w51[39] = |(datain[155:152] ^ 2);
  assign w51[40] = |(datain[151:148] ^ 3);
  assign w51[41] = |(datain[147:144] ^ 3);
  assign w51[42] = |(datain[143:140] ^ 12);
  assign w51[43] = |(datain[139:136] ^ 9);
  assign w51[44] = |(datain[135:132] ^ 9);
  assign w51[45] = |(datain[131:128] ^ 9);
  assign w51[46] = |(datain[127:124] ^ 12);
  assign w51[47] = |(datain[123:120] ^ 13);
  assign w51[48] = |(datain[119:116] ^ 2);
  assign w51[49] = |(datain[115:112] ^ 1);
  assign w51[50] = |(datain[111:108] ^ 11);
  assign w51[51] = |(datain[107:104] ^ 4);
  assign w51[52] = |(datain[103:100] ^ 2);
  assign w51[53] = |(datain[99:96] ^ 12);
  assign w51[54] = |(datain[95:92] ^ 12);
  assign w51[55] = |(datain[91:88] ^ 13);
  assign w51[56] = |(datain[87:84] ^ 2);
  assign w51[57] = |(datain[83:80] ^ 1);
  assign w51[58] = |(datain[79:76] ^ 0);
  assign w51[59] = |(datain[75:72] ^ 11);
  assign w51[60] = |(datain[71:68] ^ 13);
  assign w51[61] = |(datain[67:64] ^ 2);
  assign w51[62] = |(datain[63:60] ^ 7);
  assign w51[63] = |(datain[59:56] ^ 4);
  assign w51[64] = |(datain[55:52] ^ 15);
  assign w51[65] = |(datain[51:48] ^ 8);
  assign w51[66] = |(datain[47:44] ^ 8);
  assign w51[67] = |(datain[43:40] ^ 9);
  assign w51[68] = |(datain[39:36] ^ 9);
  assign w51[69] = |(datain[35:32] ^ 6);
  assign w51[70] = |(datain[31:28] ^ 0);
  assign w51[71] = |(datain[27:24] ^ 11);
  assign w51[72] = |(datain[23:20] ^ 0);
  assign w51[73] = |(datain[19:16] ^ 1);
  assign comp[51] = ~(|w51);
  wire [74-1:0] w52;
  assign w52[0] = |(datain[311:308] ^ 3);
  assign w52[1] = |(datain[307:304] ^ 3);
  assign w52[2] = |(datain[303:300] ^ 12);
  assign w52[3] = |(datain[299:296] ^ 9);
  assign w52[4] = |(datain[295:292] ^ 11);
  assign w52[5] = |(datain[291:288] ^ 8);
  assign w52[6] = |(datain[287:284] ^ 0);
  assign w52[7] = |(datain[283:280] ^ 0);
  assign w52[8] = |(datain[279:276] ^ 4);
  assign w52[9] = |(datain[275:272] ^ 2);
  assign w52[10] = |(datain[271:268] ^ 3);
  assign w52[11] = |(datain[267:264] ^ 3);
  assign w52[12] = |(datain[263:260] ^ 13);
  assign w52[13] = |(datain[259:256] ^ 2);
  assign w52[14] = |(datain[255:252] ^ 12);
  assign w52[15] = |(datain[251:248] ^ 13);
  assign w52[16] = |(datain[247:244] ^ 2);
  assign w52[17] = |(datain[243:240] ^ 1);
  assign w52[18] = |(datain[239:236] ^ 11);
  assign w52[19] = |(datain[235:232] ^ 10);
  assign w52[20] = |(datain[231:228] ^ 10);
  assign w52[21] = |(datain[227:224] ^ 3);
  assign w52[22] = |(datain[223:220] ^ 0);
  assign w52[23] = |(datain[219:216] ^ 4);
  assign w52[24] = |(datain[215:212] ^ 11);
  assign w52[25] = |(datain[211:208] ^ 4);
  assign w52[26] = |(datain[207:204] ^ 4);
  assign w52[27] = |(datain[203:200] ^ 0);
  assign w52[28] = |(datain[199:196] ^ 5);
  assign w52[29] = |(datain[195:192] ^ 9);
  assign w52[30] = |(datain[191:188] ^ 12);
  assign w52[31] = |(datain[187:184] ^ 13);
  assign w52[32] = |(datain[183:180] ^ 2);
  assign w52[33] = |(datain[179:176] ^ 1);
  assign w52[34] = |(datain[175:172] ^ 11);
  assign w52[35] = |(datain[171:168] ^ 8);
  assign w52[36] = |(datain[167:164] ^ 0);
  assign w52[37] = |(datain[163:160] ^ 1);
  assign w52[38] = |(datain[159:156] ^ 5);
  assign w52[39] = |(datain[155:152] ^ 7);
  assign w52[40] = |(datain[151:148] ^ 5);
  assign w52[41] = |(datain[147:144] ^ 10);
  assign w52[42] = |(datain[143:140] ^ 5);
  assign w52[43] = |(datain[139:136] ^ 9);
  assign w52[44] = |(datain[135:132] ^ 12);
  assign w52[45] = |(datain[131:128] ^ 13);
  assign w52[46] = |(datain[127:124] ^ 2);
  assign w52[47] = |(datain[123:120] ^ 1);
  assign w52[48] = |(datain[119:116] ^ 11);
  assign w52[49] = |(datain[115:112] ^ 4);
  assign w52[50] = |(datain[111:108] ^ 3);
  assign w52[51] = |(datain[107:104] ^ 14);
  assign w52[52] = |(datain[103:100] ^ 12);
  assign w52[53] = |(datain[99:96] ^ 13);
  assign w52[54] = |(datain[95:92] ^ 2);
  assign w52[55] = |(datain[91:88] ^ 1);
  assign w52[56] = |(datain[87:84] ^ 5);
  assign w52[57] = |(datain[83:80] ^ 8);
  assign w52[58] = |(datain[79:76] ^ 5);
  assign w52[59] = |(datain[75:72] ^ 10);
  assign w52[60] = |(datain[71:68] ^ 1);
  assign w52[61] = |(datain[67:64] ^ 15);
  assign w52[62] = |(datain[63:60] ^ 5);
  assign w52[63] = |(datain[59:56] ^ 9);
  assign w52[64] = |(datain[55:52] ^ 12);
  assign w52[65] = |(datain[51:48] ^ 13);
  assign w52[66] = |(datain[47:44] ^ 2);
  assign w52[67] = |(datain[43:40] ^ 1);
  assign w52[68] = |(datain[39:36] ^ 5);
  assign w52[69] = |(datain[35:32] ^ 10);
  assign w52[70] = |(datain[31:28] ^ 1);
  assign w52[71] = |(datain[27:24] ^ 15);
  assign w52[72] = |(datain[23:20] ^ 11);
  assign w52[73] = |(datain[19:16] ^ 8);
  assign comp[52] = ~(|w52);
  wire [76-1:0] w53;
  assign w53[0] = |(datain[311:308] ^ 4);
  assign w53[1] = |(datain[307:304] ^ 6);
  assign w53[2] = |(datain[303:300] ^ 14);
  assign w53[3] = |(datain[299:296] ^ 2);
  assign w53[4] = |(datain[295:292] ^ 15);
  assign w53[5] = |(datain[291:288] ^ 11);
  assign w53[6] = |(datain[287:284] ^ 11);
  assign w53[7] = |(datain[283:280] ^ 4);
  assign w53[8] = |(datain[279:276] ^ 4);
  assign w53[9] = |(datain[275:272] ^ 0);
  assign w53[10] = |(datain[271:268] ^ 11);
  assign w53[11] = |(datain[267:264] ^ 9);
  assign w53[12] = |(datain[263:260] ^ 6);
  assign w53[13] = |(datain[259:256] ^ 4);
  assign w53[14] = |(datain[255:252] ^ 0);
  assign w53[15] = |(datain[251:248] ^ 4);
  assign w53[16] = |(datain[247:244] ^ 3);
  assign w53[17] = |(datain[243:240] ^ 3);
  assign w53[18] = |(datain[239:236] ^ 13);
  assign w53[19] = |(datain[235:232] ^ 2);
  assign w53[20] = |(datain[231:228] ^ 0);
  assign w53[21] = |(datain[227:224] ^ 6);
  assign w53[22] = |(datain[223:220] ^ 1);
  assign w53[23] = |(datain[219:216] ^ 15);
  assign w53[24] = |(datain[215:212] ^ 9);
  assign w53[25] = |(datain[211:208] ^ 12);
  assign w53[26] = |(datain[207:204] ^ 2);
  assign w53[27] = |(datain[203:200] ^ 14);
  assign w53[28] = |(datain[199:196] ^ 15);
  assign w53[29] = |(datain[195:192] ^ 15);
  assign w53[30] = |(datain[191:188] ^ 1);
  assign w53[31] = |(datain[187:184] ^ 14);
  assign w53[32] = |(datain[183:180] ^ 14);
  assign w53[33] = |(datain[179:176] ^ 0);
  assign w53[34] = |(datain[175:172] ^ 0);
  assign w53[35] = |(datain[171:168] ^ 3);
  assign w53[36] = |(datain[167:164] ^ 7);
  assign w53[37] = |(datain[163:160] ^ 2);
  assign w53[38] = |(datain[159:156] ^ 3);
  assign w53[39] = |(datain[155:152] ^ 13);
  assign w53[40] = |(datain[151:148] ^ 11);
  assign w53[41] = |(datain[147:144] ^ 4);
  assign w53[42] = |(datain[143:140] ^ 4);
  assign w53[43] = |(datain[139:136] ^ 9);
  assign w53[44] = |(datain[135:132] ^ 9);
  assign w53[45] = |(datain[131:128] ^ 12);
  assign w53[46] = |(datain[127:124] ^ 2);
  assign w53[47] = |(datain[123:120] ^ 14);
  assign w53[48] = |(datain[119:116] ^ 15);
  assign w53[49] = |(datain[115:112] ^ 15);
  assign w53[50] = |(datain[111:108] ^ 1);
  assign w53[51] = |(datain[107:104] ^ 14);
  assign w53[52] = |(datain[103:100] ^ 14);
  assign w53[53] = |(datain[99:96] ^ 0);
  assign w53[54] = |(datain[95:92] ^ 0);
  assign w53[55] = |(datain[91:88] ^ 3);
  assign w53[56] = |(datain[87:84] ^ 11);
  assign w53[57] = |(datain[83:80] ^ 8);
  assign w53[58] = |(datain[79:76] ^ 0);
  assign w53[59] = |(datain[75:72] ^ 0);
  assign w53[60] = |(datain[71:68] ^ 4);
  assign w53[61] = |(datain[67:64] ^ 2);
  assign w53[62] = |(datain[63:60] ^ 9);
  assign w53[63] = |(datain[59:56] ^ 9);
  assign w53[64] = |(datain[55:52] ^ 8);
  assign w53[65] = |(datain[51:48] ^ 11);
  assign w53[66] = |(datain[47:44] ^ 12);
  assign w53[67] = |(datain[43:40] ^ 10);
  assign w53[68] = |(datain[39:36] ^ 9);
  assign w53[69] = |(datain[35:32] ^ 12);
  assign w53[70] = |(datain[31:28] ^ 2);
  assign w53[71] = |(datain[27:24] ^ 14);
  assign w53[72] = |(datain[23:20] ^ 15);
  assign w53[73] = |(datain[19:16] ^ 15);
  assign w53[74] = |(datain[15:12] ^ 1);
  assign w53[75] = |(datain[11:8] ^ 14);
  assign comp[53] = ~(|w53);
  wire [76-1:0] w54;
  assign w54[0] = |(datain[311:308] ^ 14);
  assign w54[1] = |(datain[307:304] ^ 0);
  assign w54[2] = |(datain[303:300] ^ 0);
  assign w54[3] = |(datain[299:296] ^ 3);
  assign w54[4] = |(datain[295:292] ^ 11);
  assign w54[5] = |(datain[291:288] ^ 4);
  assign w54[6] = |(datain[287:284] ^ 4);
  assign w54[7] = |(datain[283:280] ^ 0);
  assign w54[8] = |(datain[279:276] ^ 11);
  assign w54[9] = |(datain[275:272] ^ 9);
  assign w54[10] = |(datain[271:268] ^ 0);
  assign w54[11] = |(datain[267:264] ^ 3);
  assign w54[12] = |(datain[263:260] ^ 0);
  assign w54[13] = |(datain[259:256] ^ 0);
  assign w54[14] = |(datain[255:252] ^ 11);
  assign w54[15] = |(datain[251:248] ^ 10);
  assign w54[16] = |(datain[247:244] ^ 15);
  assign w54[17] = |(datain[243:240] ^ 3);
  assign w54[18] = |(datain[239:236] ^ 0);
  assign w54[19] = |(datain[235:232] ^ 3);
  assign w54[20] = |(datain[231:228] ^ 0);
  assign w54[21] = |(datain[227:224] ^ 14);
  assign w54[22] = |(datain[223:220] ^ 1);
  assign w54[23] = |(datain[219:216] ^ 15);
  assign w54[24] = |(datain[215:212] ^ 9);
  assign w54[25] = |(datain[211:208] ^ 12);
  assign w54[26] = |(datain[207:204] ^ 2);
  assign w54[27] = |(datain[203:200] ^ 14);
  assign w54[28] = |(datain[199:196] ^ 15);
  assign w54[29] = |(datain[195:192] ^ 15);
  assign w54[30] = |(datain[191:188] ^ 1);
  assign w54[31] = |(datain[187:184] ^ 14);
  assign w54[32] = |(datain[183:180] ^ 14);
  assign w54[33] = |(datain[179:176] ^ 0);
  assign w54[34] = |(datain[175:172] ^ 0);
  assign w54[35] = |(datain[171:168] ^ 3);
  assign w54[36] = |(datain[167:164] ^ 11);
  assign w54[37] = |(datain[163:160] ^ 8);
  assign w54[38] = |(datain[159:156] ^ 0);
  assign w54[39] = |(datain[155:152] ^ 1);
  assign w54[40] = |(datain[151:148] ^ 5);
  assign w54[41] = |(datain[147:144] ^ 7);
  assign w54[42] = |(datain[143:140] ^ 2);
  assign w54[43] = |(datain[139:136] ^ 14);
  assign w54[44] = |(datain[135:132] ^ 8);
  assign w54[45] = |(datain[131:128] ^ 11);
  assign w54[46] = |(datain[127:124] ^ 0);
  assign w54[47] = |(datain[123:120] ^ 14);
  assign w54[48] = |(datain[119:116] ^ 14);
  assign w54[49] = |(datain[115:112] ^ 15);
  assign w54[50] = |(datain[111:108] ^ 0);
  assign w54[51] = |(datain[107:104] ^ 3);
  assign w54[52] = |(datain[103:100] ^ 8);
  assign w54[53] = |(datain[99:96] ^ 0);
  assign w54[54] = |(datain[95:92] ^ 14);
  assign w54[55] = |(datain[91:88] ^ 1);
  assign w54[56] = |(datain[87:84] ^ 14);
  assign w54[57] = |(datain[83:80] ^ 0);
  assign w54[58] = |(datain[79:76] ^ 8);
  assign w54[59] = |(datain[75:72] ^ 0);
  assign w54[60] = |(datain[71:68] ^ 12);
  assign w54[61] = |(datain[67:64] ^ 9);
  assign w54[62] = |(datain[63:60] ^ 0);
  assign w54[63] = |(datain[59:56] ^ 13);
  assign w54[64] = |(datain[55:52] ^ 2);
  assign w54[65] = |(datain[51:48] ^ 14);
  assign w54[66] = |(datain[47:44] ^ 8);
  assign w54[67] = |(datain[43:40] ^ 11);
  assign w54[68] = |(datain[39:36] ^ 1);
  assign w54[69] = |(datain[35:32] ^ 6);
  assign w54[70] = |(datain[31:28] ^ 15);
  assign w54[71] = |(datain[27:24] ^ 1);
  assign w54[72] = |(datain[23:20] ^ 0);
  assign w54[73] = |(datain[19:16] ^ 3);
  assign w54[74] = |(datain[15:12] ^ 9);
  assign w54[75] = |(datain[11:8] ^ 12);
  assign comp[54] = ~(|w54);
  wire [74-1:0] w55;
  assign w55[0] = |(datain[311:308] ^ 14);
  assign w55[1] = |(datain[307:304] ^ 8);
  assign w55[2] = |(datain[303:300] ^ 9);
  assign w55[3] = |(datain[299:296] ^ 1);
  assign w55[4] = |(datain[295:292] ^ 0);
  assign w55[5] = |(datain[291:288] ^ 0);
  assign w55[6] = |(datain[287:284] ^ 11);
  assign w55[7] = |(datain[283:280] ^ 0);
  assign w55[8] = |(datain[279:276] ^ 0);
  assign w55[9] = |(datain[275:272] ^ 2);
  assign w55[10] = |(datain[271:268] ^ 14);
  assign w55[11] = |(datain[267:264] ^ 8);
  assign w55[12] = |(datain[263:260] ^ 8);
  assign w55[13] = |(datain[259:256] ^ 2);
  assign w55[14] = |(datain[255:252] ^ 0);
  assign w55[15] = |(datain[251:248] ^ 0);
  assign w55[16] = |(datain[247:244] ^ 11);
  assign w55[17] = |(datain[243:240] ^ 4);
  assign w55[18] = |(datain[239:236] ^ 4);
  assign w55[19] = |(datain[235:232] ^ 0);
  assign w55[20] = |(datain[231:228] ^ 8);
  assign w55[21] = |(datain[227:224] ^ 13);
  assign w55[22] = |(datain[223:220] ^ 9);
  assign w55[23] = |(datain[219:216] ^ 6);
  assign w55[24] = |(datain[215:212] ^ 7);
  assign w55[25] = |(datain[211:208] ^ 4);
  assign w55[26] = |(datain[207:204] ^ 0);
  assign w55[27] = |(datain[203:200] ^ 3);
  assign w55[28] = |(datain[199:196] ^ 5);
  assign w55[29] = |(datain[195:192] ^ 9);
  assign w55[30] = |(datain[191:188] ^ 12);
  assign w55[31] = |(datain[187:184] ^ 13);
  assign w55[32] = |(datain[183:180] ^ 2);
  assign w55[33] = |(datain[179:176] ^ 1);
  assign w55[34] = |(datain[175:172] ^ 11);
  assign w55[35] = |(datain[171:168] ^ 8);
  assign w55[36] = |(datain[167:164] ^ 0);
  assign w55[37] = |(datain[163:160] ^ 2);
  assign w55[38] = |(datain[159:156] ^ 4);
  assign w55[39] = |(datain[155:152] ^ 2);
  assign w55[40] = |(datain[151:148] ^ 3);
  assign w55[41] = |(datain[147:144] ^ 3);
  assign w55[42] = |(datain[143:140] ^ 12);
  assign w55[43] = |(datain[139:136] ^ 9);
  assign w55[44] = |(datain[135:132] ^ 9);
  assign w55[45] = |(datain[131:128] ^ 9);
  assign w55[46] = |(datain[127:124] ^ 12);
  assign w55[47] = |(datain[123:120] ^ 13);
  assign w55[48] = |(datain[119:116] ^ 2);
  assign w55[49] = |(datain[115:112] ^ 1);
  assign w55[50] = |(datain[111:108] ^ 11);
  assign w55[51] = |(datain[107:104] ^ 4);
  assign w55[52] = |(datain[103:100] ^ 2);
  assign w55[53] = |(datain[99:96] ^ 12);
  assign w55[54] = |(datain[95:92] ^ 12);
  assign w55[55] = |(datain[91:88] ^ 13);
  assign w55[56] = |(datain[87:84] ^ 2);
  assign w55[57] = |(datain[83:80] ^ 1);
  assign w55[58] = |(datain[79:76] ^ 0);
  assign w55[59] = |(datain[75:72] ^ 11);
  assign w55[60] = |(datain[71:68] ^ 13);
  assign w55[61] = |(datain[67:64] ^ 2);
  assign w55[62] = |(datain[63:60] ^ 7);
  assign w55[63] = |(datain[59:56] ^ 4);
  assign w55[64] = |(datain[55:52] ^ 15);
  assign w55[65] = |(datain[51:48] ^ 8);
  assign w55[66] = |(datain[47:44] ^ 8);
  assign w55[67] = |(datain[43:40] ^ 9);
  assign w55[68] = |(datain[39:36] ^ 9);
  assign w55[69] = |(datain[35:32] ^ 6);
  assign w55[70] = |(datain[31:28] ^ 0);
  assign w55[71] = |(datain[27:24] ^ 9);
  assign w55[72] = |(datain[23:20] ^ 0);
  assign w55[73] = |(datain[19:16] ^ 1);
  assign comp[55] = ~(|w55);
  wire [74-1:0] w56;
  assign w56[0] = |(datain[311:308] ^ 11);
  assign w56[1] = |(datain[307:304] ^ 8);
  assign w56[2] = |(datain[303:300] ^ 0);
  assign w56[3] = |(datain[299:296] ^ 0);
  assign w56[4] = |(datain[295:292] ^ 4);
  assign w56[5] = |(datain[291:288] ^ 2);
  assign w56[6] = |(datain[287:284] ^ 3);
  assign w56[7] = |(datain[283:280] ^ 3);
  assign w56[8] = |(datain[279:276] ^ 12);
  assign w56[9] = |(datain[275:272] ^ 9);
  assign w56[10] = |(datain[271:268] ^ 9);
  assign w56[11] = |(datain[267:264] ^ 9);
  assign w56[12] = |(datain[263:260] ^ 12);
  assign w56[13] = |(datain[259:256] ^ 13);
  assign w56[14] = |(datain[255:252] ^ 2);
  assign w56[15] = |(datain[251:248] ^ 1);
  assign w56[16] = |(datain[247:244] ^ 11);
  assign w56[17] = |(datain[243:240] ^ 4);
  assign w56[18] = |(datain[239:236] ^ 4);
  assign w56[19] = |(datain[235:232] ^ 0);
  assign w56[20] = |(datain[231:228] ^ 8);
  assign w56[21] = |(datain[227:224] ^ 13);
  assign w56[22] = |(datain[223:220] ^ 9);
  assign w56[23] = |(datain[219:216] ^ 6);
  assign w56[24] = |(datain[215:212] ^ 11);
  assign w56[25] = |(datain[211:208] ^ 11);
  assign w56[26] = |(datain[207:204] ^ 0);
  assign w56[27] = |(datain[203:200] ^ 2);
  assign w56[28] = |(datain[199:196] ^ 5);
  assign w56[29] = |(datain[195:192] ^ 9);
  assign w56[30] = |(datain[191:188] ^ 12);
  assign w56[31] = |(datain[187:184] ^ 13);
  assign w56[32] = |(datain[183:180] ^ 2);
  assign w56[33] = |(datain[179:176] ^ 1);
  assign w56[34] = |(datain[175:172] ^ 15);
  assign w56[35] = |(datain[171:168] ^ 14);
  assign w56[36] = |(datain[167:164] ^ 8);
  assign w56[37] = |(datain[163:160] ^ 14);
  assign w56[38] = |(datain[159:156] ^ 11);
  assign w56[39] = |(datain[155:152] ^ 10);
  assign w56[40] = |(datain[151:148] ^ 0);
  assign w56[41] = |(datain[147:144] ^ 2);
  assign w56[42] = |(datain[143:140] ^ 14);
  assign w56[43] = |(datain[139:136] ^ 9);
  assign w56[44] = |(datain[135:132] ^ 3);
  assign w56[45] = |(datain[131:128] ^ 7);
  assign w56[46] = |(datain[127:124] ^ 15);
  assign w56[47] = |(datain[123:120] ^ 15);
  assign w56[48] = |(datain[119:116] ^ 11);
  assign w56[49] = |(datain[115:112] ^ 8);
  assign w56[50] = |(datain[111:108] ^ 0);
  assign w56[51] = |(datain[107:104] ^ 1);
  assign w56[52] = |(datain[103:100] ^ 4);
  assign w56[53] = |(datain[99:96] ^ 3);
  assign w56[54] = |(datain[95:92] ^ 8);
  assign w56[55] = |(datain[91:88] ^ 13);
  assign w56[56] = |(datain[87:84] ^ 9);
  assign w56[57] = |(datain[83:80] ^ 6);
  assign w56[58] = |(datain[79:76] ^ 10);
  assign w56[59] = |(datain[75:72] ^ 13);
  assign w56[60] = |(datain[71:68] ^ 0);
  assign w56[61] = |(datain[67:64] ^ 2);
  assign w56[62] = |(datain[63:60] ^ 12);
  assign w56[63] = |(datain[59:56] ^ 13);
  assign w56[64] = |(datain[55:52] ^ 2);
  assign w56[65] = |(datain[51:48] ^ 1);
  assign w56[66] = |(datain[47:44] ^ 12);
  assign w56[67] = |(datain[43:40] ^ 3);
  assign w56[68] = |(datain[39:36] ^ 5);
  assign w56[69] = |(datain[35:32] ^ 13);
  assign w56[70] = |(datain[31:28] ^ 11);
  assign w56[71] = |(datain[27:24] ^ 4);
  assign w56[72] = |(datain[23:20] ^ 4);
  assign w56[73] = |(datain[19:16] ^ 0);
  assign comp[56] = ~(|w56);
  wire [74-1:0] w57;
  assign w57[0] = |(datain[311:308] ^ 14);
  assign w57[1] = |(datain[307:304] ^ 8);
  assign w57[2] = |(datain[303:300] ^ 8);
  assign w57[3] = |(datain[299:296] ^ 12);
  assign w57[4] = |(datain[295:292] ^ 0);
  assign w57[5] = |(datain[291:288] ^ 0);
  assign w57[6] = |(datain[287:284] ^ 11);
  assign w57[7] = |(datain[283:280] ^ 0);
  assign w57[8] = |(datain[279:276] ^ 0);
  assign w57[9] = |(datain[275:272] ^ 2);
  assign w57[10] = |(datain[271:268] ^ 14);
  assign w57[11] = |(datain[267:264] ^ 8);
  assign w57[12] = |(datain[263:260] ^ 7);
  assign w57[13] = |(datain[259:256] ^ 13);
  assign w57[14] = |(datain[255:252] ^ 0);
  assign w57[15] = |(datain[251:248] ^ 0);
  assign w57[16] = |(datain[247:244] ^ 11);
  assign w57[17] = |(datain[243:240] ^ 4);
  assign w57[18] = |(datain[239:236] ^ 4);
  assign w57[19] = |(datain[235:232] ^ 0);
  assign w57[20] = |(datain[231:228] ^ 8);
  assign w57[21] = |(datain[227:224] ^ 13);
  assign w57[22] = |(datain[223:220] ^ 9);
  assign w57[23] = |(datain[219:216] ^ 6);
  assign w57[24] = |(datain[215:212] ^ 6);
  assign w57[25] = |(datain[211:208] ^ 15);
  assign w57[26] = |(datain[207:204] ^ 0);
  assign w57[27] = |(datain[203:200] ^ 3);
  assign w57[28] = |(datain[199:196] ^ 5);
  assign w57[29] = |(datain[195:192] ^ 9);
  assign w57[30] = |(datain[191:188] ^ 12);
  assign w57[31] = |(datain[187:184] ^ 13);
  assign w57[32] = |(datain[183:180] ^ 2);
  assign w57[33] = |(datain[179:176] ^ 1);
  assign w57[34] = |(datain[175:172] ^ 11);
  assign w57[35] = |(datain[171:168] ^ 8);
  assign w57[36] = |(datain[167:164] ^ 0);
  assign w57[37] = |(datain[163:160] ^ 2);
  assign w57[38] = |(datain[159:156] ^ 4);
  assign w57[39] = |(datain[155:152] ^ 2);
  assign w57[40] = |(datain[151:148] ^ 3);
  assign w57[41] = |(datain[147:144] ^ 3);
  assign w57[42] = |(datain[143:140] ^ 12);
  assign w57[43] = |(datain[139:136] ^ 9);
  assign w57[44] = |(datain[135:132] ^ 9);
  assign w57[45] = |(datain[131:128] ^ 9);
  assign w57[46] = |(datain[127:124] ^ 12);
  assign w57[47] = |(datain[123:120] ^ 13);
  assign w57[48] = |(datain[119:116] ^ 2);
  assign w57[49] = |(datain[115:112] ^ 1);
  assign w57[50] = |(datain[111:108] ^ 11);
  assign w57[51] = |(datain[107:104] ^ 4);
  assign w57[52] = |(datain[103:100] ^ 2);
  assign w57[53] = |(datain[99:96] ^ 12);
  assign w57[54] = |(datain[95:92] ^ 12);
  assign w57[55] = |(datain[91:88] ^ 13);
  assign w57[56] = |(datain[87:84] ^ 2);
  assign w57[57] = |(datain[83:80] ^ 1);
  assign w57[58] = |(datain[79:76] ^ 0);
  assign w57[59] = |(datain[75:72] ^ 11);
  assign w57[60] = |(datain[71:68] ^ 13);
  assign w57[61] = |(datain[67:64] ^ 2);
  assign w57[62] = |(datain[63:60] ^ 7);
  assign w57[63] = |(datain[59:56] ^ 4);
  assign w57[64] = |(datain[55:52] ^ 15);
  assign w57[65] = |(datain[51:48] ^ 8);
  assign w57[66] = |(datain[47:44] ^ 8);
  assign w57[67] = |(datain[43:40] ^ 9);
  assign w57[68] = |(datain[39:36] ^ 9);
  assign w57[69] = |(datain[35:32] ^ 6);
  assign w57[70] = |(datain[31:28] ^ 0);
  assign w57[71] = |(datain[27:24] ^ 9);
  assign w57[72] = |(datain[23:20] ^ 0);
  assign w57[73] = |(datain[19:16] ^ 1);
  assign comp[57] = ~(|w57);
  wire [74-1:0] w58;
  assign w58[0] = |(datain[311:308] ^ 14);
  assign w58[1] = |(datain[307:304] ^ 8);
  assign w58[2] = |(datain[303:300] ^ 8);
  assign w58[3] = |(datain[299:296] ^ 12);
  assign w58[4] = |(datain[295:292] ^ 0);
  assign w58[5] = |(datain[291:288] ^ 0);
  assign w58[6] = |(datain[287:284] ^ 11);
  assign w58[7] = |(datain[283:280] ^ 0);
  assign w58[8] = |(datain[279:276] ^ 0);
  assign w58[9] = |(datain[275:272] ^ 2);
  assign w58[10] = |(datain[271:268] ^ 14);
  assign w58[11] = |(datain[267:264] ^ 8);
  assign w58[12] = |(datain[263:260] ^ 7);
  assign w58[13] = |(datain[259:256] ^ 13);
  assign w58[14] = |(datain[255:252] ^ 0);
  assign w58[15] = |(datain[251:248] ^ 0);
  assign w58[16] = |(datain[247:244] ^ 11);
  assign w58[17] = |(datain[243:240] ^ 4);
  assign w58[18] = |(datain[239:236] ^ 4);
  assign w58[19] = |(datain[235:232] ^ 0);
  assign w58[20] = |(datain[231:228] ^ 8);
  assign w58[21] = |(datain[227:224] ^ 13);
  assign w58[22] = |(datain[223:220] ^ 9);
  assign w58[23] = |(datain[219:216] ^ 6);
  assign w58[24] = |(datain[215:212] ^ 7);
  assign w58[25] = |(datain[211:208] ^ 2);
  assign w58[26] = |(datain[207:204] ^ 0);
  assign w58[27] = |(datain[203:200] ^ 3);
  assign w58[28] = |(datain[199:196] ^ 5);
  assign w58[29] = |(datain[195:192] ^ 9);
  assign w58[30] = |(datain[191:188] ^ 12);
  assign w58[31] = |(datain[187:184] ^ 13);
  assign w58[32] = |(datain[183:180] ^ 2);
  assign w58[33] = |(datain[179:176] ^ 1);
  assign w58[34] = |(datain[175:172] ^ 11);
  assign w58[35] = |(datain[171:168] ^ 8);
  assign w58[36] = |(datain[167:164] ^ 0);
  assign w58[37] = |(datain[163:160] ^ 2);
  assign w58[38] = |(datain[159:156] ^ 4);
  assign w58[39] = |(datain[155:152] ^ 2);
  assign w58[40] = |(datain[151:148] ^ 3);
  assign w58[41] = |(datain[147:144] ^ 3);
  assign w58[42] = |(datain[143:140] ^ 12);
  assign w58[43] = |(datain[139:136] ^ 9);
  assign w58[44] = |(datain[135:132] ^ 9);
  assign w58[45] = |(datain[131:128] ^ 9);
  assign w58[46] = |(datain[127:124] ^ 12);
  assign w58[47] = |(datain[123:120] ^ 13);
  assign w58[48] = |(datain[119:116] ^ 2);
  assign w58[49] = |(datain[115:112] ^ 1);
  assign w58[50] = |(datain[111:108] ^ 11);
  assign w58[51] = |(datain[107:104] ^ 4);
  assign w58[52] = |(datain[103:100] ^ 2);
  assign w58[53] = |(datain[99:96] ^ 12);
  assign w58[54] = |(datain[95:92] ^ 12);
  assign w58[55] = |(datain[91:88] ^ 13);
  assign w58[56] = |(datain[87:84] ^ 2);
  assign w58[57] = |(datain[83:80] ^ 1);
  assign w58[58] = |(datain[79:76] ^ 0);
  assign w58[59] = |(datain[75:72] ^ 11);
  assign w58[60] = |(datain[71:68] ^ 13);
  assign w58[61] = |(datain[67:64] ^ 2);
  assign w58[62] = |(datain[63:60] ^ 7);
  assign w58[63] = |(datain[59:56] ^ 4);
  assign w58[64] = |(datain[55:52] ^ 15);
  assign w58[65] = |(datain[51:48] ^ 8);
  assign w58[66] = |(datain[47:44] ^ 8);
  assign w58[67] = |(datain[43:40] ^ 9);
  assign w58[68] = |(datain[39:36] ^ 9);
  assign w58[69] = |(datain[35:32] ^ 6);
  assign w58[70] = |(datain[31:28] ^ 0);
  assign w58[71] = |(datain[27:24] ^ 9);
  assign w58[72] = |(datain[23:20] ^ 0);
  assign w58[73] = |(datain[19:16] ^ 1);
  assign comp[58] = ~(|w58);
  wire [76-1:0] w59;
  assign w59[0] = |(datain[311:308] ^ 11);
  assign w59[1] = |(datain[307:304] ^ 8);
  assign w59[2] = |(datain[303:300] ^ 0);
  assign w59[3] = |(datain[299:296] ^ 0);
  assign w59[4] = |(datain[295:292] ^ 4);
  assign w59[5] = |(datain[291:288] ^ 2);
  assign w59[6] = |(datain[287:284] ^ 3);
  assign w59[7] = |(datain[283:280] ^ 3);
  assign w59[8] = |(datain[279:276] ^ 12);
  assign w59[9] = |(datain[275:272] ^ 9);
  assign w59[10] = |(datain[271:268] ^ 3);
  assign w59[11] = |(datain[267:264] ^ 3);
  assign w59[12] = |(datain[263:260] ^ 13);
  assign w59[13] = |(datain[259:256] ^ 2);
  assign w59[14] = |(datain[255:252] ^ 12);
  assign w59[15] = |(datain[251:248] ^ 12);
  assign w59[16] = |(datain[247:244] ^ 8);
  assign w59[17] = |(datain[243:240] ^ 13);
  assign w59[18] = |(datain[239:236] ^ 9);
  assign w59[19] = |(datain[235:232] ^ 6);
  assign w59[20] = |(datain[231:228] ^ 4);
  assign w59[21] = |(datain[227:224] ^ 12);
  assign w59[22] = |(datain[223:220] ^ 0);
  assign w59[23] = |(datain[219:216] ^ 5);
  assign w59[24] = |(datain[215:212] ^ 11);
  assign w59[25] = |(datain[211:208] ^ 4);
  assign w59[26] = |(datain[207:204] ^ 4);
  assign w59[27] = |(datain[203:200] ^ 0);
  assign w59[28] = |(datain[199:196] ^ 11);
  assign w59[29] = |(datain[195:192] ^ 9);
  assign w59[30] = |(datain[191:188] ^ 1);
  assign w59[31] = |(datain[187:184] ^ 10);
  assign w59[32] = |(datain[183:180] ^ 0);
  assign w59[33] = |(datain[179:176] ^ 0);
  assign w59[34] = |(datain[175:172] ^ 12);
  assign w59[35] = |(datain[171:168] ^ 12);
  assign w59[36] = |(datain[167:164] ^ 15);
  assign w59[37] = |(datain[163:160] ^ 14);
  assign w59[38] = |(datain[159:156] ^ 8);
  assign w59[39] = |(datain[155:152] ^ 6);
  assign w59[40] = |(datain[151:148] ^ 4);
  assign w59[41] = |(datain[147:144] ^ 11);
  assign w59[42] = |(datain[143:140] ^ 0);
  assign w59[43] = |(datain[139:136] ^ 5);
  assign w59[44] = |(datain[135:132] ^ 11);
  assign w59[45] = |(datain[131:128] ^ 8);
  assign w59[46] = |(datain[127:124] ^ 0);
  assign w59[47] = |(datain[123:120] ^ 1);
  assign w59[48] = |(datain[119:116] ^ 5);
  assign w59[49] = |(datain[115:112] ^ 7);
  assign w59[50] = |(datain[111:108] ^ 5);
  assign w59[51] = |(datain[107:104] ^ 10);
  assign w59[52] = |(datain[103:100] ^ 5);
  assign w59[53] = |(datain[99:96] ^ 9);
  assign w59[54] = |(datain[95:92] ^ 12);
  assign w59[55] = |(datain[91:88] ^ 12);
  assign w59[56] = |(datain[87:84] ^ 11);
  assign w59[57] = |(datain[83:80] ^ 4);
  assign w59[58] = |(datain[79:76] ^ 3);
  assign w59[59] = |(datain[75:72] ^ 14);
  assign w59[60] = |(datain[71:68] ^ 12);
  assign w59[61] = |(datain[67:64] ^ 12);
  assign w59[62] = |(datain[63:60] ^ 5);
  assign w59[63] = |(datain[59:56] ^ 8);
  assign w59[64] = |(datain[55:52] ^ 5);
  assign w59[65] = |(datain[51:48] ^ 10);
  assign w59[66] = |(datain[47:44] ^ 5);
  assign w59[67] = |(datain[43:40] ^ 9);
  assign w59[68] = |(datain[39:36] ^ 12);
  assign w59[69] = |(datain[35:32] ^ 12);
  assign w59[70] = |(datain[31:28] ^ 11);
  assign w59[71] = |(datain[27:24] ^ 4);
  assign w59[72] = |(datain[23:20] ^ 4);
  assign w59[73] = |(datain[19:16] ^ 15);
  assign w59[74] = |(datain[15:12] ^ 14);
  assign w59[75] = |(datain[11:8] ^ 9);
  assign comp[59] = ~(|w59);
  wire [76-1:0] w60;
  assign w60[0] = |(datain[311:308] ^ 12);
  assign w60[1] = |(datain[307:304] ^ 9);
  assign w60[2] = |(datain[303:300] ^ 14);
  assign w60[3] = |(datain[299:296] ^ 8);
  assign w60[4] = |(datain[295:292] ^ 8);
  assign w60[5] = |(datain[291:288] ^ 12);
  assign w60[6] = |(datain[287:284] ^ 0);
  assign w60[7] = |(datain[283:280] ^ 0);
  assign w60[8] = |(datain[279:276] ^ 11);
  assign w60[9] = |(datain[275:272] ^ 0);
  assign w60[10] = |(datain[271:268] ^ 0);
  assign w60[11] = |(datain[267:264] ^ 2);
  assign w60[12] = |(datain[263:260] ^ 14);
  assign w60[13] = |(datain[259:256] ^ 8);
  assign w60[14] = |(datain[255:252] ^ 7);
  assign w60[15] = |(datain[251:248] ^ 13);
  assign w60[16] = |(datain[247:244] ^ 0);
  assign w60[17] = |(datain[243:240] ^ 0);
  assign w60[18] = |(datain[239:236] ^ 11);
  assign w60[19] = |(datain[235:232] ^ 4);
  assign w60[20] = |(datain[231:228] ^ 4);
  assign w60[21] = |(datain[227:224] ^ 0);
  assign w60[22] = |(datain[223:220] ^ 8);
  assign w60[23] = |(datain[219:216] ^ 13);
  assign w60[24] = |(datain[215:212] ^ 9);
  assign w60[25] = |(datain[211:208] ^ 6);
  assign w60[26] = |(datain[207:204] ^ 3);
  assign w60[27] = |(datain[203:200] ^ 3);
  assign w60[28] = |(datain[199:196] ^ 0);
  assign w60[29] = |(datain[195:192] ^ 4);
  assign w60[30] = |(datain[191:188] ^ 5);
  assign w60[31] = |(datain[187:184] ^ 9);
  assign w60[32] = |(datain[183:180] ^ 12);
  assign w60[33] = |(datain[179:176] ^ 13);
  assign w60[34] = |(datain[175:172] ^ 2);
  assign w60[35] = |(datain[171:168] ^ 1);
  assign w60[36] = |(datain[167:164] ^ 11);
  assign w60[37] = |(datain[163:160] ^ 8);
  assign w60[38] = |(datain[159:156] ^ 0);
  assign w60[39] = |(datain[155:152] ^ 2);
  assign w60[40] = |(datain[151:148] ^ 4);
  assign w60[41] = |(datain[147:144] ^ 2);
  assign w60[42] = |(datain[143:140] ^ 3);
  assign w60[43] = |(datain[139:136] ^ 3);
  assign w60[44] = |(datain[135:132] ^ 12);
  assign w60[45] = |(datain[131:128] ^ 9);
  assign w60[46] = |(datain[127:124] ^ 9);
  assign w60[47] = |(datain[123:120] ^ 9);
  assign w60[48] = |(datain[119:116] ^ 12);
  assign w60[49] = |(datain[115:112] ^ 13);
  assign w60[50] = |(datain[111:108] ^ 2);
  assign w60[51] = |(datain[107:104] ^ 1);
  assign w60[52] = |(datain[103:100] ^ 11);
  assign w60[53] = |(datain[99:96] ^ 4);
  assign w60[54] = |(datain[95:92] ^ 2);
  assign w60[55] = |(datain[91:88] ^ 12);
  assign w60[56] = |(datain[87:84] ^ 12);
  assign w60[57] = |(datain[83:80] ^ 13);
  assign w60[58] = |(datain[79:76] ^ 2);
  assign w60[59] = |(datain[75:72] ^ 1);
  assign w60[60] = |(datain[71:68] ^ 0);
  assign w60[61] = |(datain[67:64] ^ 11);
  assign w60[62] = |(datain[63:60] ^ 13);
  assign w60[63] = |(datain[59:56] ^ 2);
  assign w60[64] = |(datain[55:52] ^ 7);
  assign w60[65] = |(datain[51:48] ^ 4);
  assign w60[66] = |(datain[47:44] ^ 15);
  assign w60[67] = |(datain[43:40] ^ 8);
  assign w60[68] = |(datain[39:36] ^ 8);
  assign w60[69] = |(datain[35:32] ^ 9);
  assign w60[70] = |(datain[31:28] ^ 9);
  assign w60[71] = |(datain[27:24] ^ 6);
  assign w60[72] = |(datain[23:20] ^ 0);
  assign w60[73] = |(datain[19:16] ^ 11);
  assign w60[74] = |(datain[15:12] ^ 0);
  assign w60[75] = |(datain[11:8] ^ 1);
  assign comp[60] = ~(|w60);
  wire [74-1:0] w61;
  assign w61[0] = |(datain[311:308] ^ 11);
  assign w61[1] = |(datain[307:304] ^ 8);
  assign w61[2] = |(datain[303:300] ^ 0);
  assign w61[3] = |(datain[299:296] ^ 0);
  assign w61[4] = |(datain[295:292] ^ 4);
  assign w61[5] = |(datain[291:288] ^ 2);
  assign w61[6] = |(datain[287:284] ^ 3);
  assign w61[7] = |(datain[283:280] ^ 3);
  assign w61[8] = |(datain[279:276] ^ 12);
  assign w61[9] = |(datain[275:272] ^ 9);
  assign w61[10] = |(datain[271:268] ^ 9);
  assign w61[11] = |(datain[267:264] ^ 9);
  assign w61[12] = |(datain[263:260] ^ 12);
  assign w61[13] = |(datain[259:256] ^ 13);
  assign w61[14] = |(datain[255:252] ^ 2);
  assign w61[15] = |(datain[251:248] ^ 1);
  assign w61[16] = |(datain[247:244] ^ 11);
  assign w61[17] = |(datain[243:240] ^ 4);
  assign w61[18] = |(datain[239:236] ^ 4);
  assign w61[19] = |(datain[235:232] ^ 0);
  assign w61[20] = |(datain[231:228] ^ 8);
  assign w61[21] = |(datain[227:224] ^ 13);
  assign w61[22] = |(datain[223:220] ^ 9);
  assign w61[23] = |(datain[219:216] ^ 6);
  assign w61[24] = |(datain[215:212] ^ 7);
  assign w61[25] = |(datain[211:208] ^ 11);
  assign w61[26] = |(datain[207:204] ^ 0);
  assign w61[27] = |(datain[203:200] ^ 3);
  assign w61[28] = |(datain[199:196] ^ 5);
  assign w61[29] = |(datain[195:192] ^ 9);
  assign w61[30] = |(datain[191:188] ^ 12);
  assign w61[31] = |(datain[187:184] ^ 13);
  assign w61[32] = |(datain[183:180] ^ 2);
  assign w61[33] = |(datain[179:176] ^ 1);
  assign w61[34] = |(datain[175:172] ^ 15);
  assign w61[35] = |(datain[171:168] ^ 14);
  assign w61[36] = |(datain[167:164] ^ 8);
  assign w61[37] = |(datain[163:160] ^ 14);
  assign w61[38] = |(datain[159:156] ^ 7);
  assign w61[39] = |(datain[155:152] ^ 10);
  assign w61[40] = |(datain[151:148] ^ 0);
  assign w61[41] = |(datain[147:144] ^ 3);
  assign w61[42] = |(datain[143:140] ^ 14);
  assign w61[43] = |(datain[139:136] ^ 9);
  assign w61[44] = |(datain[135:132] ^ 1);
  assign w61[45] = |(datain[131:128] ^ 11);
  assign w61[46] = |(datain[127:124] ^ 15);
  assign w61[47] = |(datain[123:120] ^ 15);
  assign w61[48] = |(datain[119:116] ^ 11);
  assign w61[49] = |(datain[115:112] ^ 8);
  assign w61[50] = |(datain[111:108] ^ 0);
  assign w61[51] = |(datain[107:104] ^ 1);
  assign w61[52] = |(datain[103:100] ^ 4);
  assign w61[53] = |(datain[99:96] ^ 3);
  assign w61[54] = |(datain[95:92] ^ 8);
  assign w61[55] = |(datain[91:88] ^ 13);
  assign w61[56] = |(datain[87:84] ^ 9);
  assign w61[57] = |(datain[83:80] ^ 6);
  assign w61[58] = |(datain[79:76] ^ 6);
  assign w61[59] = |(datain[75:72] ^ 13);
  assign w61[60] = |(datain[71:68] ^ 0);
  assign w61[61] = |(datain[67:64] ^ 3);
  assign w61[62] = |(datain[63:60] ^ 12);
  assign w61[63] = |(datain[59:56] ^ 13);
  assign w61[64] = |(datain[55:52] ^ 2);
  assign w61[65] = |(datain[51:48] ^ 1);
  assign w61[66] = |(datain[47:44] ^ 12);
  assign w61[67] = |(datain[43:40] ^ 3);
  assign w61[68] = |(datain[39:36] ^ 5);
  assign w61[69] = |(datain[35:32] ^ 11);
  assign w61[70] = |(datain[31:28] ^ 11);
  assign w61[71] = |(datain[27:24] ^ 4);
  assign w61[72] = |(datain[23:20] ^ 4);
  assign w61[73] = |(datain[19:16] ^ 0);
  assign comp[61] = ~(|w61);
  wire [76-1:0] w62;
  assign w62[0] = |(datain[311:308] ^ 0);
  assign w62[1] = |(datain[307:304] ^ 6);
  assign w62[2] = |(datain[303:300] ^ 4);
  assign w62[3] = |(datain[299:296] ^ 3);
  assign w62[4] = |(datain[295:292] ^ 14);
  assign w62[5] = |(datain[291:288] ^ 8);
  assign w62[6] = |(datain[287:284] ^ 8);
  assign w62[7] = |(datain[283:280] ^ 12);
  assign w62[8] = |(datain[279:276] ^ 0);
  assign w62[9] = |(datain[275:272] ^ 1);
  assign w62[10] = |(datain[271:268] ^ 14);
  assign w62[11] = |(datain[267:264] ^ 8);
  assign w62[12] = |(datain[263:260] ^ 7);
  assign w62[13] = |(datain[259:256] ^ 5);
  assign w62[14] = |(datain[255:252] ^ 0);
  assign w62[15] = |(datain[251:248] ^ 1);
  assign w62[16] = |(datain[247:244] ^ 11);
  assign w62[17] = |(datain[243:240] ^ 4);
  assign w62[18] = |(datain[239:236] ^ 4);
  assign w62[19] = |(datain[235:232] ^ 0);
  assign w62[20] = |(datain[231:228] ^ 11);
  assign w62[21] = |(datain[227:224] ^ 9);
  assign w62[22] = |(datain[223:220] ^ 0);
  assign w62[23] = |(datain[219:216] ^ 5);
  assign w62[24] = |(datain[215:212] ^ 0);
  assign w62[25] = |(datain[211:208] ^ 0);
  assign w62[26] = |(datain[207:204] ^ 11);
  assign w62[27] = |(datain[203:200] ^ 10);
  assign w62[28] = |(datain[199:196] ^ 3);
  assign w62[29] = |(datain[195:192] ^ 4);
  assign w62[30] = |(datain[191:188] ^ 0);
  assign w62[31] = |(datain[187:184] ^ 6);
  assign w62[32] = |(datain[183:180] ^ 12);
  assign w62[33] = |(datain[179:176] ^ 13);
  assign w62[34] = |(datain[175:172] ^ 2);
  assign w62[35] = |(datain[171:168] ^ 1);
  assign w62[36] = |(datain[167:164] ^ 11);
  assign w62[37] = |(datain[163:160] ^ 8);
  assign w62[38] = |(datain[159:156] ^ 0);
  assign w62[39] = |(datain[155:152] ^ 1);
  assign w62[40] = |(datain[151:148] ^ 5);
  assign w62[41] = |(datain[147:144] ^ 7);
  assign w62[42] = |(datain[143:140] ^ 2);
  assign w62[43] = |(datain[139:136] ^ 14);
  assign w62[44] = |(datain[135:132] ^ 8);
  assign w62[45] = |(datain[131:128] ^ 11);
  assign w62[46] = |(datain[127:124] ^ 1);
  assign w62[47] = |(datain[123:120] ^ 6);
  assign w62[48] = |(datain[119:116] ^ 3);
  assign w62[49] = |(datain[115:112] ^ 11);
  assign w62[50] = |(datain[111:108] ^ 0);
  assign w62[51] = |(datain[107:104] ^ 6);
  assign w62[52] = |(datain[103:100] ^ 2);
  assign w62[53] = |(datain[99:96] ^ 14);
  assign w62[54] = |(datain[95:92] ^ 8);
  assign w62[55] = |(datain[91:88] ^ 11);
  assign w62[56] = |(datain[87:84] ^ 0);
  assign w62[57] = |(datain[83:80] ^ 14);
  assign w62[58] = |(datain[79:76] ^ 3);
  assign w62[59] = |(datain[75:72] ^ 13);
  assign w62[60] = |(datain[71:68] ^ 0);
  assign w62[61] = |(datain[67:64] ^ 6);
  assign w62[62] = |(datain[63:60] ^ 12);
  assign w62[63] = |(datain[59:56] ^ 13);
  assign w62[64] = |(datain[55:52] ^ 2);
  assign w62[65] = |(datain[51:48] ^ 1);
  assign w62[66] = |(datain[47:44] ^ 11);
  assign w62[67] = |(datain[43:40] ^ 4);
  assign w62[68] = |(datain[39:36] ^ 3);
  assign w62[69] = |(datain[35:32] ^ 14);
  assign w62[70] = |(datain[31:28] ^ 12);
  assign w62[71] = |(datain[27:24] ^ 13);
  assign w62[72] = |(datain[23:20] ^ 2);
  assign w62[73] = |(datain[19:16] ^ 1);
  assign w62[74] = |(datain[15:12] ^ 5);
  assign w62[75] = |(datain[11:8] ^ 10);
  assign comp[62] = ~(|w62);
  wire [74-1:0] w63;
  assign w63[0] = |(datain[311:308] ^ 11);
  assign w63[1] = |(datain[307:304] ^ 8);
  assign w63[2] = |(datain[303:300] ^ 0);
  assign w63[3] = |(datain[299:296] ^ 0);
  assign w63[4] = |(datain[295:292] ^ 4);
  assign w63[5] = |(datain[291:288] ^ 2);
  assign w63[6] = |(datain[287:284] ^ 3);
  assign w63[7] = |(datain[283:280] ^ 3);
  assign w63[8] = |(datain[279:276] ^ 12);
  assign w63[9] = |(datain[275:272] ^ 9);
  assign w63[10] = |(datain[271:268] ^ 9);
  assign w63[11] = |(datain[267:264] ^ 9);
  assign w63[12] = |(datain[263:260] ^ 12);
  assign w63[13] = |(datain[259:256] ^ 13);
  assign w63[14] = |(datain[255:252] ^ 2);
  assign w63[15] = |(datain[251:248] ^ 1);
  assign w63[16] = |(datain[247:244] ^ 11);
  assign w63[17] = |(datain[243:240] ^ 4);
  assign w63[18] = |(datain[239:236] ^ 4);
  assign w63[19] = |(datain[235:232] ^ 0);
  assign w63[20] = |(datain[231:228] ^ 8);
  assign w63[21] = |(datain[227:224] ^ 13);
  assign w63[22] = |(datain[223:220] ^ 9);
  assign w63[23] = |(datain[219:216] ^ 6);
  assign w63[24] = |(datain[215:212] ^ 6);
  assign w63[25] = |(datain[211:208] ^ 15);
  assign w63[26] = |(datain[207:204] ^ 0);
  assign w63[27] = |(datain[203:200] ^ 4);
  assign w63[28] = |(datain[199:196] ^ 5);
  assign w63[29] = |(datain[195:192] ^ 9);
  assign w63[30] = |(datain[191:188] ^ 12);
  assign w63[31] = |(datain[187:184] ^ 13);
  assign w63[32] = |(datain[183:180] ^ 2);
  assign w63[33] = |(datain[179:176] ^ 1);
  assign w63[34] = |(datain[175:172] ^ 15);
  assign w63[35] = |(datain[171:168] ^ 14);
  assign w63[36] = |(datain[167:164] ^ 8);
  assign w63[37] = |(datain[163:160] ^ 14);
  assign w63[38] = |(datain[159:156] ^ 6);
  assign w63[39] = |(datain[155:152] ^ 14);
  assign w63[40] = |(datain[151:148] ^ 0);
  assign w63[41] = |(datain[147:144] ^ 4);
  assign w63[42] = |(datain[143:140] ^ 14);
  assign w63[43] = |(datain[139:136] ^ 9);
  assign w63[44] = |(datain[135:132] ^ 15);
  assign w63[45] = |(datain[131:128] ^ 3);
  assign w63[46] = |(datain[127:124] ^ 15);
  assign w63[47] = |(datain[123:120] ^ 14);
  assign w63[48] = |(datain[119:116] ^ 11);
  assign w63[49] = |(datain[115:112] ^ 8);
  assign w63[50] = |(datain[111:108] ^ 0);
  assign w63[51] = |(datain[107:104] ^ 1);
  assign w63[52] = |(datain[103:100] ^ 4);
  assign w63[53] = |(datain[99:96] ^ 3);
  assign w63[54] = |(datain[95:92] ^ 8);
  assign w63[55] = |(datain[91:88] ^ 13);
  assign w63[56] = |(datain[87:84] ^ 9);
  assign w63[57] = |(datain[83:80] ^ 6);
  assign w63[58] = |(datain[79:76] ^ 6);
  assign w63[59] = |(datain[75:72] ^ 1);
  assign w63[60] = |(datain[71:68] ^ 0);
  assign w63[61] = |(datain[67:64] ^ 4);
  assign w63[62] = |(datain[63:60] ^ 12);
  assign w63[63] = |(datain[59:56] ^ 13);
  assign w63[64] = |(datain[55:52] ^ 2);
  assign w63[65] = |(datain[51:48] ^ 1);
  assign w63[66] = |(datain[47:44] ^ 12);
  assign w63[67] = |(datain[43:40] ^ 3);
  assign w63[68] = |(datain[39:36] ^ 11);
  assign w63[69] = |(datain[35:32] ^ 4);
  assign w63[70] = |(datain[31:28] ^ 4);
  assign w63[71] = |(datain[27:24] ^ 0);
  assign w63[72] = |(datain[23:20] ^ 8);
  assign w63[73] = |(datain[19:16] ^ 13);
  assign comp[63] = ~(|w63);
  wire [76-1:0] w64;
  assign w64[0] = |(datain[311:308] ^ 5);
  assign w64[1] = |(datain[307:304] ^ 7);
  assign w64[2] = |(datain[303:300] ^ 8);
  assign w64[3] = |(datain[299:296] ^ 13);
  assign w64[4] = |(datain[295:292] ^ 11);
  assign w64[5] = |(datain[291:288] ^ 6);
  assign w64[6] = |(datain[287:284] ^ 4);
  assign w64[7] = |(datain[283:280] ^ 10);
  assign w64[8] = |(datain[279:276] ^ 0);
  assign w64[9] = |(datain[275:272] ^ 1);
  assign w64[10] = |(datain[271:268] ^ 11);
  assign w64[11] = |(datain[267:264] ^ 9);
  assign w64[12] = |(datain[263:260] ^ 8);
  assign w64[13] = |(datain[259:256] ^ 10);
  assign w64[14] = |(datain[255:252] ^ 0);
  assign w64[15] = |(datain[251:248] ^ 1);
  assign w64[16] = |(datain[247:244] ^ 5);
  assign w64[17] = |(datain[243:240] ^ 1);
  assign w64[18] = |(datain[239:236] ^ 14);
  assign w64[19] = |(datain[235:232] ^ 8);
  assign w64[20] = |(datain[231:228] ^ 13);
  assign w64[21] = |(datain[227:224] ^ 5);
  assign w64[22] = |(datain[223:220] ^ 15);
  assign w64[23] = |(datain[219:216] ^ 14);
  assign w64[24] = |(datain[215:212] ^ 11);
  assign w64[25] = |(datain[211:208] ^ 4);
  assign w64[26] = |(datain[207:204] ^ 4);
  assign w64[27] = |(datain[203:200] ^ 0);
  assign w64[28] = |(datain[199:196] ^ 5);
  assign w64[29] = |(datain[195:192] ^ 9);
  assign w64[30] = |(datain[191:188] ^ 5);
  assign w64[31] = |(datain[187:184] ^ 10);
  assign w64[32] = |(datain[183:180] ^ 12);
  assign w64[33] = |(datain[179:176] ^ 13);
  assign w64[34] = |(datain[175:172] ^ 2);
  assign w64[35] = |(datain[171:168] ^ 1);
  assign w64[36] = |(datain[167:164] ^ 11);
  assign w64[37] = |(datain[163:160] ^ 8);
  assign w64[38] = |(datain[159:156] ^ 0);
  assign w64[39] = |(datain[155:152] ^ 1);
  assign w64[40] = |(datain[151:148] ^ 5);
  assign w64[41] = |(datain[147:144] ^ 7);
  assign w64[42] = |(datain[143:140] ^ 5);
  assign w64[43] = |(datain[139:136] ^ 9);
  assign w64[44] = |(datain[135:132] ^ 5);
  assign w64[45] = |(datain[131:128] ^ 10);
  assign w64[46] = |(datain[127:124] ^ 12);
  assign w64[47] = |(datain[123:120] ^ 13);
  assign w64[48] = |(datain[119:116] ^ 2);
  assign w64[49] = |(datain[115:112] ^ 1);
  assign w64[50] = |(datain[111:108] ^ 11);
  assign w64[51] = |(datain[107:104] ^ 4);
  assign w64[52] = |(datain[103:100] ^ 3);
  assign w64[53] = |(datain[99:96] ^ 14);
  assign w64[54] = |(datain[95:92] ^ 12);
  assign w64[55] = |(datain[91:88] ^ 13);
  assign w64[56] = |(datain[87:84] ^ 2);
  assign w64[57] = |(datain[83:80] ^ 1);
  assign w64[58] = |(datain[79:76] ^ 11);
  assign w64[59] = |(datain[75:72] ^ 4);
  assign w64[60] = |(datain[71:68] ^ 4);
  assign w64[61] = |(datain[67:64] ^ 15);
  assign w64[62] = |(datain[63:60] ^ 14);
  assign w64[63] = |(datain[59:56] ^ 9);
  assign w64[64] = |(datain[55:52] ^ 15);
  assign w64[65] = |(datain[51:48] ^ 13);
  assign w64[66] = |(datain[47:44] ^ 15);
  assign w64[67] = |(datain[43:40] ^ 14);
  assign w64[68] = |(datain[39:36] ^ 11);
  assign w64[69] = |(datain[35:32] ^ 8);
  assign w64[70] = |(datain[31:28] ^ 0);
  assign w64[71] = |(datain[27:24] ^ 0);
  assign w64[72] = |(datain[23:20] ^ 4);
  assign w64[73] = |(datain[19:16] ^ 2);
  assign w64[74] = |(datain[15:12] ^ 3);
  assign w64[75] = |(datain[11:8] ^ 3);
  assign comp[64] = ~(|w64);
  wire [76-1:0] w65;
  assign w65[0] = |(datain[311:308] ^ 14);
  assign w65[1] = |(datain[307:304] ^ 4);
  assign w65[2] = |(datain[303:300] ^ 4);
  assign w65[3] = |(datain[299:296] ^ 0);
  assign w65[4] = |(datain[295:292] ^ 3);
  assign w65[5] = |(datain[291:288] ^ 14);
  assign w65[6] = |(datain[287:284] ^ 8);
  assign w65[7] = |(datain[283:280] ^ 8);
  assign w65[8] = |(datain[279:276] ^ 8);
  assign w65[9] = |(datain[275:272] ^ 6);
  assign w65[10] = |(datain[271:268] ^ 4);
  assign w65[11] = |(datain[267:264] ^ 9);
  assign w65[12] = |(datain[263:260] ^ 0);
  assign w65[13] = |(datain[259:256] ^ 1);
  assign w65[14] = |(datain[255:252] ^ 11);
  assign w65[15] = |(datain[251:248] ^ 4);
  assign w65[16] = |(datain[247:244] ^ 4);
  assign w65[17] = |(datain[243:240] ^ 0);
  assign w65[18] = |(datain[239:236] ^ 8);
  assign w65[19] = |(datain[235:232] ^ 13);
  assign w65[20] = |(datain[231:228] ^ 9);
  assign w65[21] = |(datain[227:224] ^ 6);
  assign w65[22] = |(datain[223:220] ^ 0);
  assign w65[23] = |(datain[219:216] ^ 3);
  assign w65[24] = |(datain[215:212] ^ 0);
  assign w65[25] = |(datain[211:208] ^ 1);
  assign w65[26] = |(datain[207:204] ^ 11);
  assign w65[27] = |(datain[203:200] ^ 9);
  assign w65[28] = |(datain[199:196] ^ 4);
  assign w65[29] = |(datain[195:192] ^ 7);
  assign w65[30] = |(datain[191:188] ^ 0);
  assign w65[31] = |(datain[187:184] ^ 0);
  assign w65[32] = |(datain[183:180] ^ 12);
  assign w65[33] = |(datain[179:176] ^ 13);
  assign w65[34] = |(datain[175:172] ^ 2);
  assign w65[35] = |(datain[171:168] ^ 1);
  assign w65[36] = |(datain[167:164] ^ 8);
  assign w65[37] = |(datain[163:160] ^ 13);
  assign w65[38] = |(datain[159:156] ^ 11);
  assign w65[39] = |(datain[155:152] ^ 14);
  assign w65[40] = |(datain[151:148] ^ 13);
  assign w65[41] = |(datain[147:144] ^ 4);
  assign w65[42] = |(datain[143:140] ^ 0);
  assign w65[43] = |(datain[139:136] ^ 2);
  assign w65[44] = |(datain[135:132] ^ 5);
  assign w65[45] = |(datain[131:128] ^ 7);
  assign w65[46] = |(datain[127:124] ^ 8);
  assign w65[47] = |(datain[123:120] ^ 13);
  assign w65[48] = |(datain[119:116] ^ 11);
  assign w65[49] = |(datain[115:112] ^ 6);
  assign w65[50] = |(datain[111:108] ^ 4);
  assign w65[51] = |(datain[107:104] ^ 10);
  assign w65[52] = |(datain[103:100] ^ 0);
  assign w65[53] = |(datain[99:96] ^ 1);
  assign w65[54] = |(datain[95:92] ^ 11);
  assign w65[55] = |(datain[91:88] ^ 9);
  assign w65[56] = |(datain[87:84] ^ 8);
  assign w65[57] = |(datain[83:80] ^ 10);
  assign w65[58] = |(datain[79:76] ^ 0);
  assign w65[59] = |(datain[75:72] ^ 1);
  assign w65[60] = |(datain[71:68] ^ 5);
  assign w65[61] = |(datain[67:64] ^ 1);
  assign w65[62] = |(datain[63:60] ^ 14);
  assign w65[63] = |(datain[59:56] ^ 8);
  assign w65[64] = |(datain[55:52] ^ 13);
  assign w65[65] = |(datain[51:48] ^ 5);
  assign w65[66] = |(datain[47:44] ^ 15);
  assign w65[67] = |(datain[43:40] ^ 14);
  assign w65[68] = |(datain[39:36] ^ 11);
  assign w65[69] = |(datain[35:32] ^ 4);
  assign w65[70] = |(datain[31:28] ^ 4);
  assign w65[71] = |(datain[27:24] ^ 0);
  assign w65[72] = |(datain[23:20] ^ 5);
  assign w65[73] = |(datain[19:16] ^ 9);
  assign w65[74] = |(datain[15:12] ^ 5);
  assign w65[75] = |(datain[11:8] ^ 10);
  assign comp[65] = ~(|w65);
  wire [74-1:0] w66;
  assign w66[0] = |(datain[311:308] ^ 3);
  assign w66[1] = |(datain[307:304] ^ 15);
  assign w66[2] = |(datain[303:300] ^ 0);
  assign w66[3] = |(datain[299:296] ^ 3);
  assign w66[4] = |(datain[295:292] ^ 12);
  assign w66[5] = |(datain[291:288] ^ 8);
  assign w66[6] = |(datain[287:284] ^ 8);
  assign w66[7] = |(datain[283:280] ^ 9);
  assign w66[8] = |(datain[279:276] ^ 0);
  assign w66[9] = |(datain[275:272] ^ 14);
  assign w66[10] = |(datain[271:268] ^ 0);
  assign w66[11] = |(datain[267:264] ^ 4);
  assign w66[12] = |(datain[263:260] ^ 0);
  assign w66[13] = |(datain[259:256] ^ 1);
  assign w66[14] = |(datain[255:252] ^ 11);
  assign w66[15] = |(datain[251:248] ^ 4);
  assign w66[16] = |(datain[247:244] ^ 4);
  assign w66[17] = |(datain[243:240] ^ 0);
  assign w66[18] = |(datain[239:236] ^ 11);
  assign w66[19] = |(datain[235:232] ^ 10);
  assign w66[20] = |(datain[231:228] ^ 0);
  assign w66[21] = |(datain[227:224] ^ 0);
  assign w66[22] = |(datain[223:220] ^ 0);
  assign w66[23] = |(datain[219:216] ^ 1);
  assign w66[24] = |(datain[215:212] ^ 11);
  assign w66[25] = |(datain[211:208] ^ 9);
  assign w66[26] = |(datain[207:204] ^ 0);
  assign w66[27] = |(datain[203:200] ^ 12);
  assign w66[28] = |(datain[199:196] ^ 0);
  assign w66[29] = |(datain[195:192] ^ 0);
  assign w66[30] = |(datain[191:188] ^ 12);
  assign w66[31] = |(datain[187:184] ^ 13);
  assign w66[32] = |(datain[183:180] ^ 2);
  assign w66[33] = |(datain[179:176] ^ 1);
  assign w66[34] = |(datain[175:172] ^ 11);
  assign w66[35] = |(datain[171:168] ^ 4);
  assign w66[36] = |(datain[167:164] ^ 4);
  assign w66[37] = |(datain[163:160] ^ 0);
  assign w66[38] = |(datain[159:156] ^ 11);
  assign w66[39] = |(datain[155:152] ^ 10);
  assign w66[40] = |(datain[151:148] ^ 9);
  assign w66[41] = |(datain[147:144] ^ 13);
  assign w66[42] = |(datain[143:140] ^ 0);
  assign w66[43] = |(datain[139:136] ^ 1);
  assign w66[44] = |(datain[135:132] ^ 11);
  assign w66[45] = |(datain[131:128] ^ 9);
  assign w66[46] = |(datain[127:124] ^ 9);
  assign w66[47] = |(datain[123:120] ^ 1);
  assign w66[48] = |(datain[119:116] ^ 0);
  assign w66[49] = |(datain[115:112] ^ 0);
  assign w66[50] = |(datain[111:108] ^ 12);
  assign w66[51] = |(datain[107:104] ^ 13);
  assign w66[52] = |(datain[103:100] ^ 2);
  assign w66[53] = |(datain[99:96] ^ 1);
  assign w66[54] = |(datain[95:92] ^ 11);
  assign w66[55] = |(datain[91:88] ^ 4);
  assign w66[56] = |(datain[87:84] ^ 3);
  assign w66[57] = |(datain[83:80] ^ 14);
  assign w66[58] = |(datain[79:76] ^ 12);
  assign w66[59] = |(datain[75:72] ^ 13);
  assign w66[60] = |(datain[71:68] ^ 2);
  assign w66[61] = |(datain[67:64] ^ 1);
  assign w66[62] = |(datain[63:60] ^ 11);
  assign w66[63] = |(datain[59:56] ^ 4);
  assign w66[64] = |(datain[55:52] ^ 4);
  assign w66[65] = |(datain[51:48] ^ 15);
  assign w66[66] = |(datain[47:44] ^ 14);
  assign w66[67] = |(datain[43:40] ^ 11);
  assign w66[68] = |(datain[39:36] ^ 8);
  assign w66[69] = |(datain[35:32] ^ 6);
  assign w66[70] = |(datain[31:28] ^ 11);
  assign w66[71] = |(datain[27:24] ^ 4);
  assign w66[72] = |(datain[23:20] ^ 0);
  assign w66[73] = |(datain[19:16] ^ 9);
  assign comp[66] = ~(|w66);
  wire [76-1:0] w67;
  assign w67[0] = |(datain[311:308] ^ 5);
  assign w67[1] = |(datain[307:304] ^ 11);
  assign w67[2] = |(datain[303:300] ^ 11);
  assign w67[3] = |(datain[299:296] ^ 4);
  assign w67[4] = |(datain[295:292] ^ 4);
  assign w67[5] = |(datain[291:288] ^ 0);
  assign w67[6] = |(datain[287:284] ^ 11);
  assign w67[7] = |(datain[283:280] ^ 9);
  assign w67[8] = |(datain[279:276] ^ 3);
  assign w67[9] = |(datain[275:272] ^ 15);
  assign w67[10] = |(datain[271:268] ^ 0);
  assign w67[11] = |(datain[267:264] ^ 4);
  assign w67[12] = |(datain[263:260] ^ 11);
  assign w67[13] = |(datain[259:256] ^ 10);
  assign w67[14] = |(datain[255:252] ^ 4);
  assign w67[15] = |(datain[251:248] ^ 6);
  assign w67[16] = |(datain[247:244] ^ 0);
  assign w67[17] = |(datain[243:240] ^ 5);
  assign w67[18] = |(datain[239:236] ^ 12);
  assign w67[19] = |(datain[235:232] ^ 13);
  assign w67[20] = |(datain[231:228] ^ 0);
  assign w67[21] = |(datain[227:224] ^ 1);
  assign w67[22] = |(datain[223:220] ^ 11);
  assign w67[23] = |(datain[219:216] ^ 8);
  assign w67[24] = |(datain[215:212] ^ 0);
  assign w67[25] = |(datain[211:208] ^ 0);
  assign w67[26] = |(datain[207:204] ^ 4);
  assign w67[27] = |(datain[203:200] ^ 2);
  assign w67[28] = |(datain[199:196] ^ 3);
  assign w67[29] = |(datain[195:192] ^ 3);
  assign w67[30] = |(datain[191:188] ^ 12);
  assign w67[31] = |(datain[187:184] ^ 9);
  assign w67[32] = |(datain[183:180] ^ 3);
  assign w67[33] = |(datain[179:176] ^ 3);
  assign w67[34] = |(datain[175:172] ^ 13);
  assign w67[35] = |(datain[171:168] ^ 2);
  assign w67[36] = |(datain[167:164] ^ 12);
  assign w67[37] = |(datain[163:160] ^ 13);
  assign w67[38] = |(datain[159:156] ^ 0);
  assign w67[39] = |(datain[155:152] ^ 1);
  assign w67[40] = |(datain[151:148] ^ 11);
  assign w67[41] = |(datain[147:144] ^ 4);
  assign w67[42] = |(datain[143:140] ^ 4);
  assign w67[43] = |(datain[139:136] ^ 0);
  assign w67[44] = |(datain[135:132] ^ 11);
  assign w67[45] = |(datain[131:128] ^ 10);
  assign w67[46] = |(datain[127:124] ^ 4);
  assign w67[47] = |(datain[123:120] ^ 3);
  assign w67[48] = |(datain[119:116] ^ 0);
  assign w67[49] = |(datain[115:112] ^ 5);
  assign w67[50] = |(datain[111:108] ^ 11);
  assign w67[51] = |(datain[107:104] ^ 9);
  assign w67[52] = |(datain[103:100] ^ 0);
  assign w67[53] = |(datain[99:96] ^ 3);
  assign w67[54] = |(datain[95:92] ^ 0);
  assign w67[55] = |(datain[91:88] ^ 0);
  assign w67[56] = |(datain[87:84] ^ 12);
  assign w67[57] = |(datain[83:80] ^ 12);
  assign w67[58] = |(datain[79:76] ^ 5);
  assign w67[59] = |(datain[75:72] ^ 10);
  assign w67[60] = |(datain[71:68] ^ 5);
  assign w67[61] = |(datain[67:64] ^ 9);
  assign w67[62] = |(datain[63:60] ^ 11);
  assign w67[63] = |(datain[59:56] ^ 8);
  assign w67[64] = |(datain[55:52] ^ 0);
  assign w67[65] = |(datain[51:48] ^ 1);
  assign w67[66] = |(datain[47:44] ^ 5);
  assign w67[67] = |(datain[43:40] ^ 7);
  assign w67[68] = |(datain[39:36] ^ 12);
  assign w67[69] = |(datain[35:32] ^ 13);
  assign w67[70] = |(datain[31:28] ^ 0);
  assign w67[71] = |(datain[27:24] ^ 1);
  assign w67[72] = |(datain[23:20] ^ 11);
  assign w67[73] = |(datain[19:16] ^ 4);
  assign w67[74] = |(datain[15:12] ^ 3);
  assign w67[75] = |(datain[11:8] ^ 14);
  assign comp[67] = ~(|w67);
  wire [74-1:0] w68;
  assign w68[0] = |(datain[311:308] ^ 14);
  assign w68[1] = |(datain[307:304] ^ 8);
  assign w68[2] = |(datain[303:300] ^ 8);
  assign w68[3] = |(datain[299:296] ^ 12);
  assign w68[4] = |(datain[295:292] ^ 0);
  assign w68[5] = |(datain[291:288] ^ 0);
  assign w68[6] = |(datain[287:284] ^ 11);
  assign w68[7] = |(datain[283:280] ^ 0);
  assign w68[8] = |(datain[279:276] ^ 0);
  assign w68[9] = |(datain[275:272] ^ 2);
  assign w68[10] = |(datain[271:268] ^ 14);
  assign w68[11] = |(datain[267:264] ^ 8);
  assign w68[12] = |(datain[263:260] ^ 7);
  assign w68[13] = |(datain[259:256] ^ 13);
  assign w68[14] = |(datain[255:252] ^ 0);
  assign w68[15] = |(datain[251:248] ^ 0);
  assign w68[16] = |(datain[247:244] ^ 11);
  assign w68[17] = |(datain[243:240] ^ 4);
  assign w68[18] = |(datain[239:236] ^ 4);
  assign w68[19] = |(datain[235:232] ^ 0);
  assign w68[20] = |(datain[231:228] ^ 8);
  assign w68[21] = |(datain[227:224] ^ 13);
  assign w68[22] = |(datain[223:220] ^ 9);
  assign w68[23] = |(datain[219:216] ^ 6);
  assign w68[24] = |(datain[215:212] ^ 7);
  assign w68[25] = |(datain[211:208] ^ 5);
  assign w68[26] = |(datain[207:204] ^ 0);
  assign w68[27] = |(datain[203:200] ^ 3);
  assign w68[28] = |(datain[199:196] ^ 5);
  assign w68[29] = |(datain[195:192] ^ 9);
  assign w68[30] = |(datain[191:188] ^ 12);
  assign w68[31] = |(datain[187:184] ^ 13);
  assign w68[32] = |(datain[183:180] ^ 2);
  assign w68[33] = |(datain[179:176] ^ 1);
  assign w68[34] = |(datain[175:172] ^ 11);
  assign w68[35] = |(datain[171:168] ^ 8);
  assign w68[36] = |(datain[167:164] ^ 0);
  assign w68[37] = |(datain[163:160] ^ 2);
  assign w68[38] = |(datain[159:156] ^ 4);
  assign w68[39] = |(datain[155:152] ^ 2);
  assign w68[40] = |(datain[151:148] ^ 3);
  assign w68[41] = |(datain[147:144] ^ 3);
  assign w68[42] = |(datain[143:140] ^ 12);
  assign w68[43] = |(datain[139:136] ^ 9);
  assign w68[44] = |(datain[135:132] ^ 9);
  assign w68[45] = |(datain[131:128] ^ 9);
  assign w68[46] = |(datain[127:124] ^ 12);
  assign w68[47] = |(datain[123:120] ^ 13);
  assign w68[48] = |(datain[119:116] ^ 2);
  assign w68[49] = |(datain[115:112] ^ 1);
  assign w68[50] = |(datain[111:108] ^ 11);
  assign w68[51] = |(datain[107:104] ^ 4);
  assign w68[52] = |(datain[103:100] ^ 2);
  assign w68[53] = |(datain[99:96] ^ 12);
  assign w68[54] = |(datain[95:92] ^ 12);
  assign w68[55] = |(datain[91:88] ^ 13);
  assign w68[56] = |(datain[87:84] ^ 2);
  assign w68[57] = |(datain[83:80] ^ 1);
  assign w68[58] = |(datain[79:76] ^ 0);
  assign w68[59] = |(datain[75:72] ^ 11);
  assign w68[60] = |(datain[71:68] ^ 13);
  assign w68[61] = |(datain[67:64] ^ 2);
  assign w68[62] = |(datain[63:60] ^ 7);
  assign w68[63] = |(datain[59:56] ^ 4);
  assign w68[64] = |(datain[55:52] ^ 15);
  assign w68[65] = |(datain[51:48] ^ 8);
  assign w68[66] = |(datain[47:44] ^ 8);
  assign w68[67] = |(datain[43:40] ^ 9);
  assign w68[68] = |(datain[39:36] ^ 9);
  assign w68[69] = |(datain[35:32] ^ 6);
  assign w68[70] = |(datain[31:28] ^ 0);
  assign w68[71] = |(datain[27:24] ^ 10);
  assign w68[72] = |(datain[23:20] ^ 0);
  assign w68[73] = |(datain[19:16] ^ 1);
  assign comp[68] = ~(|w68);
  wire [74-1:0] w69;
  assign w69[0] = |(datain[311:308] ^ 14);
  assign w69[1] = |(datain[307:304] ^ 8);
  assign w69[2] = |(datain[303:300] ^ 8);
  assign w69[3] = |(datain[299:296] ^ 12);
  assign w69[4] = |(datain[295:292] ^ 0);
  assign w69[5] = |(datain[291:288] ^ 0);
  assign w69[6] = |(datain[287:284] ^ 11);
  assign w69[7] = |(datain[283:280] ^ 0);
  assign w69[8] = |(datain[279:276] ^ 0);
  assign w69[9] = |(datain[275:272] ^ 2);
  assign w69[10] = |(datain[271:268] ^ 14);
  assign w69[11] = |(datain[267:264] ^ 8);
  assign w69[12] = |(datain[263:260] ^ 7);
  assign w69[13] = |(datain[259:256] ^ 13);
  assign w69[14] = |(datain[255:252] ^ 0);
  assign w69[15] = |(datain[251:248] ^ 0);
  assign w69[16] = |(datain[247:244] ^ 11);
  assign w69[17] = |(datain[243:240] ^ 4);
  assign w69[18] = |(datain[239:236] ^ 4);
  assign w69[19] = |(datain[235:232] ^ 0);
  assign w69[20] = |(datain[231:228] ^ 8);
  assign w69[21] = |(datain[227:224] ^ 13);
  assign w69[22] = |(datain[223:220] ^ 9);
  assign w69[23] = |(datain[219:216] ^ 6);
  assign w69[24] = |(datain[215:212] ^ 8);
  assign w69[25] = |(datain[211:208] ^ 2);
  assign w69[26] = |(datain[207:204] ^ 0);
  assign w69[27] = |(datain[203:200] ^ 3);
  assign w69[28] = |(datain[199:196] ^ 5);
  assign w69[29] = |(datain[195:192] ^ 9);
  assign w69[30] = |(datain[191:188] ^ 12);
  assign w69[31] = |(datain[187:184] ^ 13);
  assign w69[32] = |(datain[183:180] ^ 2);
  assign w69[33] = |(datain[179:176] ^ 1);
  assign w69[34] = |(datain[175:172] ^ 11);
  assign w69[35] = |(datain[171:168] ^ 8);
  assign w69[36] = |(datain[167:164] ^ 0);
  assign w69[37] = |(datain[163:160] ^ 2);
  assign w69[38] = |(datain[159:156] ^ 4);
  assign w69[39] = |(datain[155:152] ^ 2);
  assign w69[40] = |(datain[151:148] ^ 3);
  assign w69[41] = |(datain[147:144] ^ 3);
  assign w69[42] = |(datain[143:140] ^ 12);
  assign w69[43] = |(datain[139:136] ^ 9);
  assign w69[44] = |(datain[135:132] ^ 9);
  assign w69[45] = |(datain[131:128] ^ 9);
  assign w69[46] = |(datain[127:124] ^ 12);
  assign w69[47] = |(datain[123:120] ^ 13);
  assign w69[48] = |(datain[119:116] ^ 2);
  assign w69[49] = |(datain[115:112] ^ 1);
  assign w69[50] = |(datain[111:108] ^ 11);
  assign w69[51] = |(datain[107:104] ^ 4);
  assign w69[52] = |(datain[103:100] ^ 2);
  assign w69[53] = |(datain[99:96] ^ 12);
  assign w69[54] = |(datain[95:92] ^ 12);
  assign w69[55] = |(datain[91:88] ^ 13);
  assign w69[56] = |(datain[87:84] ^ 2);
  assign w69[57] = |(datain[83:80] ^ 1);
  assign w69[58] = |(datain[79:76] ^ 0);
  assign w69[59] = |(datain[75:72] ^ 11);
  assign w69[60] = |(datain[71:68] ^ 13);
  assign w69[61] = |(datain[67:64] ^ 2);
  assign w69[62] = |(datain[63:60] ^ 7);
  assign w69[63] = |(datain[59:56] ^ 4);
  assign w69[64] = |(datain[55:52] ^ 15);
  assign w69[65] = |(datain[51:48] ^ 8);
  assign w69[66] = |(datain[47:44] ^ 8);
  assign w69[67] = |(datain[43:40] ^ 9);
  assign w69[68] = |(datain[39:36] ^ 9);
  assign w69[69] = |(datain[35:32] ^ 6);
  assign w69[70] = |(datain[31:28] ^ 0);
  assign w69[71] = |(datain[27:24] ^ 11);
  assign w69[72] = |(datain[23:20] ^ 0);
  assign w69[73] = |(datain[19:16] ^ 1);
  assign comp[69] = ~(|w69);
  wire [76-1:0] w70;
  assign w70[0] = |(datain[311:308] ^ 10);
  assign w70[1] = |(datain[307:304] ^ 3);
  assign w70[2] = |(datain[303:300] ^ 0);
  assign w70[3] = |(datain[299:296] ^ 6);
  assign w70[4] = |(datain[295:292] ^ 0);
  assign w70[5] = |(datain[291:288] ^ 1);
  assign w70[6] = |(datain[287:284] ^ 11);
  assign w70[7] = |(datain[283:280] ^ 4);
  assign w70[8] = |(datain[279:276] ^ 4);
  assign w70[9] = |(datain[275:272] ^ 0);
  assign w70[10] = |(datain[271:268] ^ 12);
  assign w70[11] = |(datain[267:264] ^ 13);
  assign w70[12] = |(datain[263:260] ^ 2);
  assign w70[13] = |(datain[259:256] ^ 1);
  assign w70[14] = |(datain[255:252] ^ 3);
  assign w70[15] = |(datain[251:248] ^ 2);
  assign w70[16] = |(datain[247:244] ^ 12);
  assign w70[17] = |(datain[243:240] ^ 0);
  assign w70[18] = |(datain[239:236] ^ 14);
  assign w70[19] = |(datain[235:232] ^ 8);
  assign w70[20] = |(datain[231:228] ^ 1);
  assign w70[21] = |(datain[227:224] ^ 2);
  assign w70[22] = |(datain[223:220] ^ 0);
  assign w70[23] = |(datain[219:216] ^ 0);
  assign w70[24] = |(datain[215:212] ^ 8);
  assign w70[25] = |(datain[211:208] ^ 11);
  assign w70[26] = |(datain[207:204] ^ 13);
  assign w70[27] = |(datain[203:200] ^ 7);
  assign w70[28] = |(datain[199:196] ^ 11);
  assign w70[29] = |(datain[195:192] ^ 4);
  assign w70[30] = |(datain[191:188] ^ 4);
  assign w70[31] = |(datain[187:184] ^ 0);
  assign w70[32] = |(datain[183:180] ^ 12);
  assign w70[33] = |(datain[179:176] ^ 13);
  assign w70[34] = |(datain[175:172] ^ 2);
  assign w70[35] = |(datain[171:168] ^ 1);
  assign w70[36] = |(datain[167:164] ^ 11);
  assign w70[37] = |(datain[163:160] ^ 4);
  assign w70[38] = |(datain[159:156] ^ 3);
  assign w70[39] = |(datain[155:152] ^ 14);
  assign w70[40] = |(datain[151:148] ^ 12);
  assign w70[41] = |(datain[147:144] ^ 13);
  assign w70[42] = |(datain[143:140] ^ 2);
  assign w70[43] = |(datain[139:136] ^ 1);
  assign w70[44] = |(datain[135:132] ^ 11);
  assign w70[45] = |(datain[131:128] ^ 4);
  assign w70[46] = |(datain[127:124] ^ 4);
  assign w70[47] = |(datain[123:120] ^ 15);
  assign w70[48] = |(datain[119:116] ^ 14);
  assign w70[49] = |(datain[115:112] ^ 11);
  assign w70[50] = |(datain[111:108] ^ 12);
  assign w70[51] = |(datain[107:104] ^ 7);
  assign w70[52] = |(datain[103:100] ^ 5);
  assign w70[53] = |(datain[99:96] ^ 7);
  assign w70[54] = |(datain[95:92] ^ 15);
  assign w70[55] = |(datain[91:88] ^ 3);
  assign w70[56] = |(datain[87:84] ^ 10);
  assign w70[57] = |(datain[83:80] ^ 4);
  assign w70[58] = |(datain[79:76] ^ 12);
  assign w70[59] = |(datain[75:72] ^ 3);
  assign w70[60] = |(datain[71:68] ^ 5);
  assign w70[61] = |(datain[67:64] ^ 1);
  assign w70[62] = |(datain[63:60] ^ 5);
  assign w70[63] = |(datain[59:56] ^ 2);
  assign w70[64] = |(datain[55:52] ^ 9);
  assign w70[65] = |(datain[51:48] ^ 9);
  assign w70[66] = |(datain[47:44] ^ 3);
  assign w70[67] = |(datain[43:40] ^ 3);
  assign w70[68] = |(datain[39:36] ^ 12);
  assign w70[69] = |(datain[35:32] ^ 9);
  assign w70[70] = |(datain[31:28] ^ 11);
  assign w70[71] = |(datain[27:24] ^ 4);
  assign w70[72] = |(datain[23:20] ^ 4);
  assign w70[73] = |(datain[19:16] ^ 2);
  assign w70[74] = |(datain[15:12] ^ 12);
  assign w70[75] = |(datain[11:8] ^ 13);
  assign comp[70] = ~(|w70);
  wire [76-1:0] w71;
  assign w71[0] = |(datain[311:308] ^ 12);
  assign w71[1] = |(datain[307:304] ^ 9);
  assign w71[2] = |(datain[303:300] ^ 14);
  assign w71[3] = |(datain[299:296] ^ 8);
  assign w71[4] = |(datain[295:292] ^ 9);
  assign w71[5] = |(datain[291:288] ^ 1);
  assign w71[6] = |(datain[287:284] ^ 0);
  assign w71[7] = |(datain[283:280] ^ 0);
  assign w71[8] = |(datain[279:276] ^ 11);
  assign w71[9] = |(datain[275:272] ^ 0);
  assign w71[10] = |(datain[271:268] ^ 0);
  assign w71[11] = |(datain[267:264] ^ 2);
  assign w71[12] = |(datain[263:260] ^ 14);
  assign w71[13] = |(datain[259:256] ^ 8);
  assign w71[14] = |(datain[255:252] ^ 8);
  assign w71[15] = |(datain[251:248] ^ 2);
  assign w71[16] = |(datain[247:244] ^ 0);
  assign w71[17] = |(datain[243:240] ^ 0);
  assign w71[18] = |(datain[239:236] ^ 11);
  assign w71[19] = |(datain[235:232] ^ 4);
  assign w71[20] = |(datain[231:228] ^ 4);
  assign w71[21] = |(datain[227:224] ^ 0);
  assign w71[22] = |(datain[223:220] ^ 8);
  assign w71[23] = |(datain[219:216] ^ 13);
  assign w71[24] = |(datain[215:212] ^ 9);
  assign w71[25] = |(datain[211:208] ^ 6);
  assign w71[26] = |(datain[207:204] ^ 7);
  assign w71[27] = |(datain[203:200] ^ 10);
  assign w71[28] = |(datain[199:196] ^ 0);
  assign w71[29] = |(datain[195:192] ^ 3);
  assign w71[30] = |(datain[191:188] ^ 5);
  assign w71[31] = |(datain[187:184] ^ 9);
  assign w71[32] = |(datain[183:180] ^ 12);
  assign w71[33] = |(datain[179:176] ^ 13);
  assign w71[34] = |(datain[175:172] ^ 2);
  assign w71[35] = |(datain[171:168] ^ 1);
  assign w71[36] = |(datain[167:164] ^ 11);
  assign w71[37] = |(datain[163:160] ^ 8);
  assign w71[38] = |(datain[159:156] ^ 0);
  assign w71[39] = |(datain[155:152] ^ 2);
  assign w71[40] = |(datain[151:148] ^ 4);
  assign w71[41] = |(datain[147:144] ^ 2);
  assign w71[42] = |(datain[143:140] ^ 3);
  assign w71[43] = |(datain[139:136] ^ 3);
  assign w71[44] = |(datain[135:132] ^ 12);
  assign w71[45] = |(datain[131:128] ^ 9);
  assign w71[46] = |(datain[127:124] ^ 9);
  assign w71[47] = |(datain[123:120] ^ 9);
  assign w71[48] = |(datain[119:116] ^ 12);
  assign w71[49] = |(datain[115:112] ^ 13);
  assign w71[50] = |(datain[111:108] ^ 2);
  assign w71[51] = |(datain[107:104] ^ 1);
  assign w71[52] = |(datain[103:100] ^ 11);
  assign w71[53] = |(datain[99:96] ^ 4);
  assign w71[54] = |(datain[95:92] ^ 2);
  assign w71[55] = |(datain[91:88] ^ 12);
  assign w71[56] = |(datain[87:84] ^ 12);
  assign w71[57] = |(datain[83:80] ^ 13);
  assign w71[58] = |(datain[79:76] ^ 2);
  assign w71[59] = |(datain[75:72] ^ 1);
  assign w71[60] = |(datain[71:68] ^ 0);
  assign w71[61] = |(datain[67:64] ^ 11);
  assign w71[62] = |(datain[63:60] ^ 13);
  assign w71[63] = |(datain[59:56] ^ 2);
  assign w71[64] = |(datain[55:52] ^ 7);
  assign w71[65] = |(datain[51:48] ^ 4);
  assign w71[66] = |(datain[47:44] ^ 15);
  assign w71[67] = |(datain[43:40] ^ 8);
  assign w71[68] = |(datain[39:36] ^ 8);
  assign w71[69] = |(datain[35:32] ^ 9);
  assign w71[70] = |(datain[31:28] ^ 9);
  assign w71[71] = |(datain[27:24] ^ 6);
  assign w71[72] = |(datain[23:20] ^ 0);
  assign w71[73] = |(datain[19:16] ^ 10);
  assign w71[74] = |(datain[15:12] ^ 0);
  assign w71[75] = |(datain[11:8] ^ 1);
  assign comp[71] = ~(|w71);
  wire [74-1:0] w72;
  assign w72[0] = |(datain[311:308] ^ 14);
  assign w72[1] = |(datain[307:304] ^ 8);
  assign w72[2] = |(datain[303:300] ^ 11);
  assign w72[3] = |(datain[299:296] ^ 13);
  assign w72[4] = |(datain[295:292] ^ 15);
  assign w72[5] = |(datain[291:288] ^ 15);
  assign w72[6] = |(datain[287:284] ^ 11);
  assign w72[7] = |(datain[283:280] ^ 0);
  assign w72[8] = |(datain[279:276] ^ 0);
  assign w72[9] = |(datain[275:272] ^ 2);
  assign w72[10] = |(datain[271:268] ^ 14);
  assign w72[11] = |(datain[267:264] ^ 8);
  assign w72[12] = |(datain[263:260] ^ 7);
  assign w72[13] = |(datain[259:256] ^ 8);
  assign w72[14] = |(datain[255:252] ^ 15);
  assign w72[15] = |(datain[251:248] ^ 15);
  assign w72[16] = |(datain[247:244] ^ 11);
  assign w72[17] = |(datain[243:240] ^ 4);
  assign w72[18] = |(datain[239:236] ^ 4);
  assign w72[19] = |(datain[235:232] ^ 0);
  assign w72[20] = |(datain[231:228] ^ 8);
  assign w72[21] = |(datain[227:224] ^ 13);
  assign w72[22] = |(datain[223:220] ^ 9);
  assign w72[23] = |(datain[219:216] ^ 6);
  assign w72[24] = |(datain[215:212] ^ 10);
  assign w72[25] = |(datain[211:208] ^ 11);
  assign w72[26] = |(datain[207:204] ^ 0);
  assign w72[27] = |(datain[203:200] ^ 2);
  assign w72[28] = |(datain[199:196] ^ 5);
  assign w72[29] = |(datain[195:192] ^ 9);
  assign w72[30] = |(datain[191:188] ^ 12);
  assign w72[31] = |(datain[187:184] ^ 13);
  assign w72[32] = |(datain[183:180] ^ 2);
  assign w72[33] = |(datain[179:176] ^ 1);
  assign w72[34] = |(datain[175:172] ^ 11);
  assign w72[35] = |(datain[171:168] ^ 8);
  assign w72[36] = |(datain[167:164] ^ 0);
  assign w72[37] = |(datain[163:160] ^ 2);
  assign w72[38] = |(datain[159:156] ^ 4);
  assign w72[39] = |(datain[155:152] ^ 2);
  assign w72[40] = |(datain[151:148] ^ 3);
  assign w72[41] = |(datain[147:144] ^ 3);
  assign w72[42] = |(datain[143:140] ^ 12);
  assign w72[43] = |(datain[139:136] ^ 9);
  assign w72[44] = |(datain[135:132] ^ 9);
  assign w72[45] = |(datain[131:128] ^ 9);
  assign w72[46] = |(datain[127:124] ^ 12);
  assign w72[47] = |(datain[123:120] ^ 13);
  assign w72[48] = |(datain[119:116] ^ 2);
  assign w72[49] = |(datain[115:112] ^ 1);
  assign w72[50] = |(datain[111:108] ^ 11);
  assign w72[51] = |(datain[107:104] ^ 4);
  assign w72[52] = |(datain[103:100] ^ 2);
  assign w72[53] = |(datain[99:96] ^ 12);
  assign w72[54] = |(datain[95:92] ^ 12);
  assign w72[55] = |(datain[91:88] ^ 13);
  assign w72[56] = |(datain[87:84] ^ 2);
  assign w72[57] = |(datain[83:80] ^ 1);
  assign w72[58] = |(datain[79:76] ^ 0);
  assign w72[59] = |(datain[75:72] ^ 11);
  assign w72[60] = |(datain[71:68] ^ 13);
  assign w72[61] = |(datain[67:64] ^ 2);
  assign w72[62] = |(datain[63:60] ^ 7);
  assign w72[63] = |(datain[59:56] ^ 4);
  assign w72[64] = |(datain[55:52] ^ 15);
  assign w72[65] = |(datain[51:48] ^ 8);
  assign w72[66] = |(datain[47:44] ^ 8);
  assign w72[67] = |(datain[43:40] ^ 9);
  assign w72[68] = |(datain[39:36] ^ 8);
  assign w72[69] = |(datain[35:32] ^ 14);
  assign w72[70] = |(datain[31:28] ^ 0);
  assign w72[71] = |(datain[27:24] ^ 11);
  assign w72[72] = |(datain[23:20] ^ 0);
  assign w72[73] = |(datain[19:16] ^ 1);
  assign comp[72] = ~(|w72);
  wire [74-1:0] w73;
  assign w73[0] = |(datain[311:308] ^ 11);
  assign w73[1] = |(datain[307:304] ^ 14);
  assign w73[2] = |(datain[303:300] ^ 0);
  assign w73[3] = |(datain[299:296] ^ 5);
  assign w73[4] = |(datain[295:292] ^ 0);
  assign w73[5] = |(datain[291:288] ^ 1);
  assign w73[6] = |(datain[287:284] ^ 11);
  assign w73[7] = |(datain[283:280] ^ 9);
  assign w73[8] = |(datain[279:276] ^ 11);
  assign w73[9] = |(datain[275:272] ^ 3);
  assign w73[10] = |(datain[271:268] ^ 0);
  assign w73[11] = |(datain[267:264] ^ 6);
  assign w73[12] = |(datain[263:260] ^ 9);
  assign w73[13] = |(datain[259:256] ^ 0);
  assign w73[14] = |(datain[255:252] ^ 0);
  assign w73[15] = |(datain[251:248] ^ 5);
  assign w73[16] = |(datain[247:244] ^ 0);
  assign w73[17] = |(datain[243:240] ^ 3);
  assign w73[18] = |(datain[239:236] ^ 0);
  assign w73[19] = |(datain[235:232] ^ 1);
  assign w73[20] = |(datain[231:228] ^ 8);
  assign w73[21] = |(datain[227:224] ^ 11);
  assign w73[22] = |(datain[223:220] ^ 13);
  assign w73[23] = |(datain[219:216] ^ 0);
  assign w73[24] = |(datain[215:212] ^ 14);
  assign w73[25] = |(datain[211:208] ^ 8);
  assign w73[26] = |(datain[207:204] ^ 5);
  assign w73[27] = |(datain[203:200] ^ 1);
  assign w73[28] = |(datain[199:196] ^ 0);
  assign w73[29] = |(datain[195:192] ^ 0);
  assign w73[30] = |(datain[191:188] ^ 5);
  assign w73[31] = |(datain[187:184] ^ 15);
  assign w73[32] = |(datain[183:180] ^ 0);
  assign w73[33] = |(datain[179:176] ^ 7);
  assign w73[34] = |(datain[175:172] ^ 11);
  assign w73[35] = |(datain[171:168] ^ 4);
  assign w73[36] = |(datain[167:164] ^ 4);
  assign w73[37] = |(datain[163:160] ^ 0);
  assign w73[38] = |(datain[159:156] ^ 12);
  assign w73[39] = |(datain[155:152] ^ 13);
  assign w73[40] = |(datain[151:148] ^ 2);
  assign w73[41] = |(datain[147:144] ^ 1);
  assign w73[42] = |(datain[143:140] ^ 2);
  assign w73[43] = |(datain[139:136] ^ 6);
  assign w73[44] = |(datain[135:132] ^ 12);
  assign w73[45] = |(datain[131:128] ^ 7);
  assign w73[46] = |(datain[127:124] ^ 4);
  assign w73[47] = |(datain[123:120] ^ 5);
  assign w73[48] = |(datain[119:116] ^ 1);
  assign w73[49] = |(datain[115:112] ^ 5);
  assign w73[50] = |(datain[111:108] ^ 0);
  assign w73[51] = |(datain[107:104] ^ 0);
  assign w73[52] = |(datain[103:100] ^ 0);
  assign w73[53] = |(datain[99:96] ^ 0);
  assign w73[54] = |(datain[95:92] ^ 11);
  assign w73[55] = |(datain[91:88] ^ 4);
  assign w73[56] = |(datain[87:84] ^ 4);
  assign w73[57] = |(datain[83:80] ^ 0);
  assign w73[58] = |(datain[79:76] ^ 11);
  assign w73[59] = |(datain[75:72] ^ 10);
  assign w73[60] = |(datain[71:68] ^ 4);
  assign w73[61] = |(datain[67:64] ^ 9);
  assign w73[62] = |(datain[63:60] ^ 0);
  assign w73[63] = |(datain[59:56] ^ 2);
  assign w73[64] = |(datain[55:52] ^ 11);
  assign w73[65] = |(datain[51:48] ^ 9);
  assign w73[66] = |(datain[47:44] ^ 0);
  assign w73[67] = |(datain[43:40] ^ 5);
  assign w73[68] = |(datain[39:36] ^ 0);
  assign w73[69] = |(datain[35:32] ^ 0);
  assign w73[70] = |(datain[31:28] ^ 12);
  assign w73[71] = |(datain[27:24] ^ 13);
  assign w73[72] = |(datain[23:20] ^ 2);
  assign w73[73] = |(datain[19:16] ^ 1);
  assign comp[73] = ~(|w73);
  wire [74-1:0] w74;
  assign w74[0] = |(datain[311:308] ^ 12);
  assign w74[1] = |(datain[307:304] ^ 13);
  assign w74[2] = |(datain[303:300] ^ 2);
  assign w74[3] = |(datain[299:296] ^ 1);
  assign w74[4] = |(datain[295:292] ^ 11);
  assign w74[5] = |(datain[291:288] ^ 4);
  assign w74[6] = |(datain[287:284] ^ 4);
  assign w74[7] = |(datain[283:280] ^ 0);
  assign w74[8] = |(datain[279:276] ^ 2);
  assign w74[9] = |(datain[275:272] ^ 14);
  assign w74[10] = |(datain[271:268] ^ 8);
  assign w74[11] = |(datain[267:264] ^ 11);
  assign w74[12] = |(datain[263:260] ^ 1);
  assign w74[13] = |(datain[259:256] ^ 14);
  assign w74[14] = |(datain[255:252] ^ 1);
  assign w74[15] = |(datain[251:248] ^ 13);
  assign w74[16] = |(datain[247:244] ^ 0);
  assign w74[17] = |(datain[243:240] ^ 1);
  assign w74[18] = |(datain[239:236] ^ 11);
  assign w74[19] = |(datain[235:232] ^ 9);
  assign w74[20] = |(datain[231:228] ^ 12);
  assign w74[21] = |(datain[227:224] ^ 12);
  assign w74[22] = |(datain[223:220] ^ 0);
  assign w74[23] = |(datain[219:216] ^ 1);
  assign w74[24] = |(datain[215:212] ^ 11);
  assign w74[25] = |(datain[211:208] ^ 10);
  assign w74[26] = |(datain[207:204] ^ 0);
  assign w74[27] = |(datain[203:200] ^ 0);
  assign w74[28] = |(datain[199:196] ^ 0);
  assign w74[29] = |(datain[195:192] ^ 1);
  assign w74[30] = |(datain[191:188] ^ 12);
  assign w74[31] = |(datain[187:184] ^ 13);
  assign w74[32] = |(datain[183:180] ^ 2);
  assign w74[33] = |(datain[179:176] ^ 1);
  assign w74[34] = |(datain[175:172] ^ 11);
  assign w74[35] = |(datain[171:168] ^ 8);
  assign w74[36] = |(datain[167:164] ^ 0);
  assign w74[37] = |(datain[163:160] ^ 0);
  assign w74[38] = |(datain[159:156] ^ 4);
  assign w74[39] = |(datain[155:152] ^ 2);
  assign w74[40] = |(datain[151:148] ^ 2);
  assign w74[41] = |(datain[147:144] ^ 14);
  assign w74[42] = |(datain[143:140] ^ 8);
  assign w74[43] = |(datain[139:136] ^ 11);
  assign w74[44] = |(datain[135:132] ^ 1);
  assign w74[45] = |(datain[131:128] ^ 14);
  assign w74[46] = |(datain[127:124] ^ 1);
  assign w74[47] = |(datain[123:120] ^ 13);
  assign w74[48] = |(datain[119:116] ^ 0);
  assign w74[49] = |(datain[115:112] ^ 1);
  assign w74[50] = |(datain[111:108] ^ 3);
  assign w74[51] = |(datain[107:104] ^ 3);
  assign w74[52] = |(datain[103:100] ^ 12);
  assign w74[53] = |(datain[99:96] ^ 9);
  assign w74[54] = |(datain[95:92] ^ 3);
  assign w74[55] = |(datain[91:88] ^ 3);
  assign w74[56] = |(datain[87:84] ^ 13);
  assign w74[57] = |(datain[83:80] ^ 2);
  assign w74[58] = |(datain[79:76] ^ 12);
  assign w74[59] = |(datain[75:72] ^ 13);
  assign w74[60] = |(datain[71:68] ^ 2);
  assign w74[61] = |(datain[67:64] ^ 1);
  assign w74[62] = |(datain[63:60] ^ 2);
  assign w74[63] = |(datain[59:56] ^ 14);
  assign w74[64] = |(datain[55:52] ^ 10);
  assign w74[65] = |(datain[51:48] ^ 1);
  assign w74[66] = |(datain[47:44] ^ 1);
  assign w74[67] = |(datain[43:40] ^ 15);
  assign w74[68] = |(datain[39:36] ^ 0);
  assign w74[69] = |(datain[35:32] ^ 1);
  assign w74[70] = |(datain[31:28] ^ 2);
  assign w74[71] = |(datain[27:24] ^ 13);
  assign w74[72] = |(datain[23:20] ^ 0);
  assign w74[73] = |(datain[19:16] ^ 3);
  assign comp[74] = ~(|w74);
  wire [74-1:0] w75;
  assign w75[0] = |(datain[311:308] ^ 2);
  assign w75[1] = |(datain[307:304] ^ 14);
  assign w75[2] = |(datain[303:300] ^ 2);
  assign w75[3] = |(datain[299:296] ^ 11);
  assign w75[4] = |(datain[295:292] ^ 0);
  assign w75[5] = |(datain[291:288] ^ 14);
  assign w75[6] = |(datain[287:284] ^ 1);
  assign w75[7] = |(datain[283:280] ^ 15);
  assign w75[8] = |(datain[279:276] ^ 0);
  assign w75[9] = |(datain[275:272] ^ 1);
  assign w75[10] = |(datain[271:268] ^ 11);
  assign w75[11] = |(datain[267:264] ^ 4);
  assign w75[12] = |(datain[263:260] ^ 4);
  assign w75[13] = |(datain[259:256] ^ 0);
  assign w75[14] = |(datain[255:252] ^ 2);
  assign w75[15] = |(datain[251:248] ^ 14);
  assign w75[16] = |(datain[247:244] ^ 8);
  assign w75[17] = |(datain[243:240] ^ 11);
  assign w75[18] = |(datain[239:236] ^ 1);
  assign w75[19] = |(datain[235:232] ^ 14);
  assign w75[20] = |(datain[231:228] ^ 1);
  assign w75[21] = |(datain[227:224] ^ 13);
  assign w75[22] = |(datain[223:220] ^ 0);
  assign w75[23] = |(datain[219:216] ^ 1);
  assign w75[24] = |(datain[215:212] ^ 11);
  assign w75[25] = |(datain[211:208] ^ 10);
  assign w75[26] = |(datain[207:204] ^ 4);
  assign w75[27] = |(datain[203:200] ^ 7);
  assign w75[28] = |(datain[199:196] ^ 0);
  assign w75[29] = |(datain[195:192] ^ 1);
  assign w75[30] = |(datain[191:188] ^ 12);
  assign w75[31] = |(datain[187:184] ^ 13);
  assign w75[32] = |(datain[183:180] ^ 2);
  assign w75[33] = |(datain[179:176] ^ 1);
  assign w75[34] = |(datain[175:172] ^ 11);
  assign w75[35] = |(datain[171:168] ^ 4);
  assign w75[36] = |(datain[167:164] ^ 4);
  assign w75[37] = |(datain[163:160] ^ 0);
  assign w75[38] = |(datain[159:156] ^ 2);
  assign w75[39] = |(datain[155:152] ^ 14);
  assign w75[40] = |(datain[151:148] ^ 8);
  assign w75[41] = |(datain[147:144] ^ 11);
  assign w75[42] = |(datain[143:140] ^ 1);
  assign w75[43] = |(datain[139:136] ^ 14);
  assign w75[44] = |(datain[135:132] ^ 1);
  assign w75[45] = |(datain[131:128] ^ 13);
  assign w75[46] = |(datain[127:124] ^ 0);
  assign w75[47] = |(datain[123:120] ^ 1);
  assign w75[48] = |(datain[119:116] ^ 11);
  assign w75[49] = |(datain[115:112] ^ 9);
  assign w75[50] = |(datain[111:108] ^ 12);
  assign w75[51] = |(datain[107:104] ^ 12);
  assign w75[52] = |(datain[103:100] ^ 0);
  assign w75[53] = |(datain[99:96] ^ 1);
  assign w75[54] = |(datain[95:92] ^ 11);
  assign w75[55] = |(datain[91:88] ^ 10);
  assign w75[56] = |(datain[87:84] ^ 0);
  assign w75[57] = |(datain[83:80] ^ 0);
  assign w75[58] = |(datain[79:76] ^ 0);
  assign w75[59] = |(datain[75:72] ^ 1);
  assign w75[60] = |(datain[71:68] ^ 12);
  assign w75[61] = |(datain[67:64] ^ 13);
  assign w75[62] = |(datain[63:60] ^ 2);
  assign w75[63] = |(datain[59:56] ^ 1);
  assign w75[64] = |(datain[55:52] ^ 11);
  assign w75[65] = |(datain[51:48] ^ 8);
  assign w75[66] = |(datain[47:44] ^ 0);
  assign w75[67] = |(datain[43:40] ^ 0);
  assign w75[68] = |(datain[39:36] ^ 4);
  assign w75[69] = |(datain[35:32] ^ 2);
  assign w75[70] = |(datain[31:28] ^ 2);
  assign w75[71] = |(datain[27:24] ^ 14);
  assign w75[72] = |(datain[23:20] ^ 8);
  assign w75[73] = |(datain[19:16] ^ 11);
  assign comp[75] = ~(|w75);
  wire [76-1:0] w76;
  assign w76[0] = |(datain[311:308] ^ 0);
  assign w76[1] = |(datain[307:304] ^ 8);
  assign w76[2] = |(datain[303:300] ^ 11);
  assign w76[3] = |(datain[299:296] ^ 14);
  assign w76[4] = |(datain[295:292] ^ 0);
  assign w76[5] = |(datain[291:288] ^ 5);
  assign w76[6] = |(datain[287:284] ^ 0);
  assign w76[7] = |(datain[283:280] ^ 1);
  assign w76[8] = |(datain[279:276] ^ 11);
  assign w76[9] = |(datain[275:272] ^ 9);
  assign w76[10] = |(datain[271:268] ^ 11);
  assign w76[11] = |(datain[267:264] ^ 14);
  assign w76[12] = |(datain[263:260] ^ 0);
  assign w76[13] = |(datain[259:256] ^ 7);
  assign w76[14] = |(datain[255:252] ^ 9);
  assign w76[15] = |(datain[251:248] ^ 0);
  assign w76[16] = |(datain[247:244] ^ 0);
  assign w76[17] = |(datain[243:240] ^ 5);
  assign w76[18] = |(datain[239:236] ^ 0);
  assign w76[19] = |(datain[235:232] ^ 3);
  assign w76[20] = |(datain[231:228] ^ 0);
  assign w76[21] = |(datain[227:224] ^ 1);
  assign w76[22] = |(datain[223:220] ^ 8);
  assign w76[23] = |(datain[219:216] ^ 11);
  assign w76[24] = |(datain[215:212] ^ 13);
  assign w76[25] = |(datain[211:208] ^ 0);
  assign w76[26] = |(datain[207:204] ^ 14);
  assign w76[27] = |(datain[203:200] ^ 8);
  assign w76[28] = |(datain[199:196] ^ 5);
  assign w76[29] = |(datain[195:192] ^ 1);
  assign w76[30] = |(datain[191:188] ^ 0);
  assign w76[31] = |(datain[187:184] ^ 0);
  assign w76[32] = |(datain[183:180] ^ 5);
  assign w76[33] = |(datain[179:176] ^ 15);
  assign w76[34] = |(datain[175:172] ^ 0);
  assign w76[35] = |(datain[171:168] ^ 7);
  assign w76[36] = |(datain[167:164] ^ 11);
  assign w76[37] = |(datain[163:160] ^ 4);
  assign w76[38] = |(datain[159:156] ^ 4);
  assign w76[39] = |(datain[155:152] ^ 0);
  assign w76[40] = |(datain[151:148] ^ 12);
  assign w76[41] = |(datain[147:144] ^ 13);
  assign w76[42] = |(datain[143:140] ^ 2);
  assign w76[43] = |(datain[139:136] ^ 1);
  assign w76[44] = |(datain[135:132] ^ 2);
  assign w76[45] = |(datain[131:128] ^ 6);
  assign w76[46] = |(datain[127:124] ^ 12);
  assign w76[47] = |(datain[123:120] ^ 7);
  assign w76[48] = |(datain[119:116] ^ 4);
  assign w76[49] = |(datain[115:112] ^ 5);
  assign w76[50] = |(datain[111:108] ^ 1);
  assign w76[51] = |(datain[107:104] ^ 5);
  assign w76[52] = |(datain[103:100] ^ 0);
  assign w76[53] = |(datain[99:96] ^ 0);
  assign w76[54] = |(datain[95:92] ^ 0);
  assign w76[55] = |(datain[91:88] ^ 0);
  assign w76[56] = |(datain[87:84] ^ 11);
  assign w76[57] = |(datain[83:80] ^ 4);
  assign w76[58] = |(datain[79:76] ^ 4);
  assign w76[59] = |(datain[75:72] ^ 0);
  assign w76[60] = |(datain[71:68] ^ 11);
  assign w76[61] = |(datain[67:64] ^ 10);
  assign w76[62] = |(datain[63:60] ^ 4);
  assign w76[63] = |(datain[59:56] ^ 9);
  assign w76[64] = |(datain[55:52] ^ 0);
  assign w76[65] = |(datain[51:48] ^ 2);
  assign w76[66] = |(datain[47:44] ^ 11);
  assign w76[67] = |(datain[43:40] ^ 9);
  assign w76[68] = |(datain[39:36] ^ 0);
  assign w76[69] = |(datain[35:32] ^ 5);
  assign w76[70] = |(datain[31:28] ^ 0);
  assign w76[71] = |(datain[27:24] ^ 0);
  assign w76[72] = |(datain[23:20] ^ 12);
  assign w76[73] = |(datain[19:16] ^ 13);
  assign w76[74] = |(datain[15:12] ^ 2);
  assign w76[75] = |(datain[11:8] ^ 1);
  assign comp[76] = ~(|w76);
  wire [76-1:0] w77;
  assign w77[0] = |(datain[311:308] ^ 0);
  assign w77[1] = |(datain[307:304] ^ 8);
  assign w77[2] = |(datain[303:300] ^ 11);
  assign w77[3] = |(datain[299:296] ^ 14);
  assign w77[4] = |(datain[295:292] ^ 0);
  assign w77[5] = |(datain[291:288] ^ 5);
  assign w77[6] = |(datain[287:284] ^ 0);
  assign w77[7] = |(datain[283:280] ^ 1);
  assign w77[8] = |(datain[279:276] ^ 11);
  assign w77[9] = |(datain[275:272] ^ 9);
  assign w77[10] = |(datain[271:268] ^ 5);
  assign w77[11] = |(datain[267:264] ^ 2);
  assign w77[12] = |(datain[263:260] ^ 0);
  assign w77[13] = |(datain[259:256] ^ 7);
  assign w77[14] = |(datain[255:252] ^ 9);
  assign w77[15] = |(datain[251:248] ^ 0);
  assign w77[16] = |(datain[247:244] ^ 0);
  assign w77[17] = |(datain[243:240] ^ 5);
  assign w77[18] = |(datain[239:236] ^ 0);
  assign w77[19] = |(datain[235:232] ^ 3);
  assign w77[20] = |(datain[231:228] ^ 0);
  assign w77[21] = |(datain[227:224] ^ 1);
  assign w77[22] = |(datain[223:220] ^ 8);
  assign w77[23] = |(datain[219:216] ^ 11);
  assign w77[24] = |(datain[215:212] ^ 13);
  assign w77[25] = |(datain[211:208] ^ 0);
  assign w77[26] = |(datain[207:204] ^ 14);
  assign w77[27] = |(datain[203:200] ^ 8);
  assign w77[28] = |(datain[199:196] ^ 5);
  assign w77[29] = |(datain[195:192] ^ 1);
  assign w77[30] = |(datain[191:188] ^ 0);
  assign w77[31] = |(datain[187:184] ^ 0);
  assign w77[32] = |(datain[183:180] ^ 5);
  assign w77[33] = |(datain[179:176] ^ 15);
  assign w77[34] = |(datain[175:172] ^ 0);
  assign w77[35] = |(datain[171:168] ^ 7);
  assign w77[36] = |(datain[167:164] ^ 11);
  assign w77[37] = |(datain[163:160] ^ 4);
  assign w77[38] = |(datain[159:156] ^ 4);
  assign w77[39] = |(datain[155:152] ^ 0);
  assign w77[40] = |(datain[151:148] ^ 12);
  assign w77[41] = |(datain[147:144] ^ 13);
  assign w77[42] = |(datain[143:140] ^ 2);
  assign w77[43] = |(datain[139:136] ^ 1);
  assign w77[44] = |(datain[135:132] ^ 2);
  assign w77[45] = |(datain[131:128] ^ 6);
  assign w77[46] = |(datain[127:124] ^ 12);
  assign w77[47] = |(datain[123:120] ^ 7);
  assign w77[48] = |(datain[119:116] ^ 4);
  assign w77[49] = |(datain[115:112] ^ 5);
  assign w77[50] = |(datain[111:108] ^ 1);
  assign w77[51] = |(datain[107:104] ^ 5);
  assign w77[52] = |(datain[103:100] ^ 0);
  assign w77[53] = |(datain[99:96] ^ 0);
  assign w77[54] = |(datain[95:92] ^ 0);
  assign w77[55] = |(datain[91:88] ^ 0);
  assign w77[56] = |(datain[87:84] ^ 11);
  assign w77[57] = |(datain[83:80] ^ 4);
  assign w77[58] = |(datain[79:76] ^ 4);
  assign w77[59] = |(datain[75:72] ^ 0);
  assign w77[60] = |(datain[71:68] ^ 11);
  assign w77[61] = |(datain[67:64] ^ 10);
  assign w77[62] = |(datain[63:60] ^ 4);
  assign w77[63] = |(datain[59:56] ^ 9);
  assign w77[64] = |(datain[55:52] ^ 0);
  assign w77[65] = |(datain[51:48] ^ 2);
  assign w77[66] = |(datain[47:44] ^ 11);
  assign w77[67] = |(datain[43:40] ^ 9);
  assign w77[68] = |(datain[39:36] ^ 0);
  assign w77[69] = |(datain[35:32] ^ 5);
  assign w77[70] = |(datain[31:28] ^ 0);
  assign w77[71] = |(datain[27:24] ^ 0);
  assign w77[72] = |(datain[23:20] ^ 12);
  assign w77[73] = |(datain[19:16] ^ 13);
  assign w77[74] = |(datain[15:12] ^ 2);
  assign w77[75] = |(datain[11:8] ^ 1);
  assign comp[77] = ~(|w77);
  wire [74-1:0] w78;
  assign w78[0] = |(datain[311:308] ^ 3);
  assign w78[1] = |(datain[307:304] ^ 3);
  assign w78[2] = |(datain[303:300] ^ 12);
  assign w78[3] = |(datain[299:296] ^ 9);
  assign w78[4] = |(datain[295:292] ^ 3);
  assign w78[5] = |(datain[291:288] ^ 3);
  assign w78[6] = |(datain[287:284] ^ 13);
  assign w78[7] = |(datain[283:280] ^ 2);
  assign w78[8] = |(datain[279:276] ^ 12);
  assign w78[9] = |(datain[275:272] ^ 13);
  assign w78[10] = |(datain[271:268] ^ 2);
  assign w78[11] = |(datain[267:264] ^ 1);
  assign w78[12] = |(datain[263:260] ^ 11);
  assign w78[13] = |(datain[259:256] ^ 4);
  assign w78[14] = |(datain[255:252] ^ 4);
  assign w78[15] = |(datain[251:248] ^ 0);
  assign w78[16] = |(datain[247:244] ^ 11);
  assign w78[17] = |(datain[243:240] ^ 9);
  assign w78[18] = |(datain[239:236] ^ 7);
  assign w78[19] = |(datain[235:232] ^ 2);
  assign w78[20] = |(datain[231:228] ^ 0);
  assign w78[21] = |(datain[227:224] ^ 1);
  assign w78[22] = |(datain[223:220] ^ 8);
  assign w78[23] = |(datain[219:216] ^ 13);
  assign w78[24] = |(datain[215:212] ^ 9);
  assign w78[25] = |(datain[211:208] ^ 6);
  assign w78[26] = |(datain[207:204] ^ 0);
  assign w78[27] = |(datain[203:200] ^ 5);
  assign w78[28] = |(datain[199:196] ^ 0);
  assign w78[29] = |(datain[195:192] ^ 0);
  assign w78[30] = |(datain[191:188] ^ 12);
  assign w78[31] = |(datain[187:184] ^ 13);
  assign w78[32] = |(datain[183:180] ^ 2);
  assign w78[33] = |(datain[179:176] ^ 1);
  assign w78[34] = |(datain[175:172] ^ 14);
  assign w78[35] = |(datain[171:168] ^ 8);
  assign w78[36] = |(datain[167:164] ^ 2);
  assign w78[37] = |(datain[163:160] ^ 8);
  assign w78[38] = |(datain[159:156] ^ 0);
  assign w78[39] = |(datain[155:152] ^ 0);
  assign w78[40] = |(datain[151:148] ^ 8);
  assign w78[41] = |(datain[147:144] ^ 13);
  assign w78[42] = |(datain[143:140] ^ 9);
  assign w78[43] = |(datain[139:136] ^ 6);
  assign w78[44] = |(datain[135:132] ^ 9);
  assign w78[45] = |(datain[131:128] ^ 1);
  assign w78[46] = |(datain[127:124] ^ 0);
  assign w78[47] = |(datain[123:120] ^ 1);
  assign w78[48] = |(datain[119:116] ^ 11);
  assign w78[49] = |(datain[115:112] ^ 4);
  assign w78[50] = |(datain[111:108] ^ 0);
  assign w78[51] = |(datain[107:104] ^ 9);
  assign w78[52] = |(datain[103:100] ^ 12);
  assign w78[53] = |(datain[99:96] ^ 13);
  assign w78[54] = |(datain[95:92] ^ 2);
  assign w78[55] = |(datain[91:88] ^ 1);
  assign w78[56] = |(datain[87:84] ^ 8);
  assign w78[57] = |(datain[83:80] ^ 13);
  assign w78[58] = |(datain[79:76] ^ 9);
  assign w78[59] = |(datain[75:72] ^ 6);
  assign w78[60] = |(datain[71:68] ^ 7);
  assign w78[61] = |(datain[67:64] ^ 0);
  assign w78[62] = |(datain[63:60] ^ 0);
  assign w78[63] = |(datain[59:56] ^ 1);
  assign w78[64] = |(datain[55:52] ^ 12);
  assign w78[65] = |(datain[51:48] ^ 13);
  assign w78[66] = |(datain[47:44] ^ 2);
  assign w78[67] = |(datain[43:40] ^ 1);
  assign w78[68] = |(datain[39:36] ^ 12);
  assign w78[69] = |(datain[35:32] ^ 3);
  assign w78[70] = |(datain[31:28] ^ 11);
  assign w78[71] = |(datain[27:24] ^ 9);
  assign w78[72] = |(datain[23:20] ^ 2);
  assign w78[73] = |(datain[19:16] ^ 0);
  assign comp[78] = ~(|w78);
  wire [76-1:0] w79;
  assign w79[0] = |(datain[311:308] ^ 4);
  assign w79[1] = |(datain[307:304] ^ 2);
  assign w79[2] = |(datain[303:300] ^ 3);
  assign w79[3] = |(datain[299:296] ^ 3);
  assign w79[4] = |(datain[295:292] ^ 12);
  assign w79[5] = |(datain[291:288] ^ 9);
  assign w79[6] = |(datain[287:284] ^ 3);
  assign w79[7] = |(datain[283:280] ^ 3);
  assign w79[8] = |(datain[279:276] ^ 13);
  assign w79[9] = |(datain[275:272] ^ 2);
  assign w79[10] = |(datain[271:268] ^ 12);
  assign w79[11] = |(datain[267:264] ^ 13);
  assign w79[12] = |(datain[263:260] ^ 2);
  assign w79[13] = |(datain[259:256] ^ 1);
  assign w79[14] = |(datain[255:252] ^ 11);
  assign w79[15] = |(datain[251:248] ^ 4);
  assign w79[16] = |(datain[247:244] ^ 4);
  assign w79[17] = |(datain[243:240] ^ 0);
  assign w79[18] = |(datain[239:236] ^ 11);
  assign w79[19] = |(datain[235:232] ^ 9);
  assign w79[20] = |(datain[231:228] ^ 0);
  assign w79[21] = |(datain[227:224] ^ 5);
  assign w79[22] = |(datain[223:220] ^ 0);
  assign w79[23] = |(datain[219:216] ^ 0);
  assign w79[24] = |(datain[215:212] ^ 8);
  assign w79[25] = |(datain[211:208] ^ 13);
  assign w79[26] = |(datain[207:204] ^ 9);
  assign w79[27] = |(datain[203:200] ^ 6);
  assign w79[28] = |(datain[199:196] ^ 11);
  assign w79[29] = |(datain[195:192] ^ 3);
  assign w79[30] = |(datain[191:188] ^ 0);
  assign w79[31] = |(datain[187:184] ^ 0);
  assign w79[32] = |(datain[183:180] ^ 12);
  assign w79[33] = |(datain[179:176] ^ 13);
  assign w79[34] = |(datain[175:172] ^ 2);
  assign w79[35] = |(datain[171:168] ^ 1);
  assign w79[36] = |(datain[167:164] ^ 11);
  assign w79[37] = |(datain[163:160] ^ 8);
  assign w79[38] = |(datain[159:156] ^ 0);
  assign w79[39] = |(datain[155:152] ^ 2);
  assign w79[40] = |(datain[151:148] ^ 4);
  assign w79[41] = |(datain[147:144] ^ 2);
  assign w79[42] = |(datain[143:140] ^ 3);
  assign w79[43] = |(datain[139:136] ^ 3);
  assign w79[44] = |(datain[135:132] ^ 12);
  assign w79[45] = |(datain[131:128] ^ 9);
  assign w79[46] = |(datain[127:124] ^ 3);
  assign w79[47] = |(datain[123:120] ^ 3);
  assign w79[48] = |(datain[119:116] ^ 13);
  assign w79[49] = |(datain[115:112] ^ 2);
  assign w79[50] = |(datain[111:108] ^ 12);
  assign w79[51] = |(datain[107:104] ^ 13);
  assign w79[52] = |(datain[103:100] ^ 2);
  assign w79[53] = |(datain[99:96] ^ 1);
  assign w79[54] = |(datain[95:92] ^ 11);
  assign w79[55] = |(datain[91:88] ^ 4);
  assign w79[56] = |(datain[87:84] ^ 4);
  assign w79[57] = |(datain[83:80] ^ 0);
  assign w79[58] = |(datain[79:76] ^ 11);
  assign w79[59] = |(datain[75:72] ^ 9);
  assign w79[60] = |(datain[71:68] ^ 7);
  assign w79[61] = |(datain[67:64] ^ 2);
  assign w79[62] = |(datain[63:60] ^ 0);
  assign w79[63] = |(datain[59:56] ^ 1);
  assign w79[64] = |(datain[55:52] ^ 8);
  assign w79[65] = |(datain[51:48] ^ 13);
  assign w79[66] = |(datain[47:44] ^ 9);
  assign w79[67] = |(datain[43:40] ^ 6);
  assign w79[68] = |(datain[39:36] ^ 0);
  assign w79[69] = |(datain[35:32] ^ 5);
  assign w79[70] = |(datain[31:28] ^ 0);
  assign w79[71] = |(datain[27:24] ^ 0);
  assign w79[72] = |(datain[23:20] ^ 12);
  assign w79[73] = |(datain[19:16] ^ 13);
  assign w79[74] = |(datain[15:12] ^ 2);
  assign w79[75] = |(datain[11:8] ^ 1);
  assign comp[79] = ~(|w79);
  wire [74-1:0] w80;
  assign w80[0] = |(datain[311:308] ^ 4);
  assign w80[1] = |(datain[307:304] ^ 2);
  assign w80[2] = |(datain[303:300] ^ 3);
  assign w80[3] = |(datain[299:296] ^ 3);
  assign w80[4] = |(datain[295:292] ^ 12);
  assign w80[5] = |(datain[291:288] ^ 9);
  assign w80[6] = |(datain[287:284] ^ 3);
  assign w80[7] = |(datain[283:280] ^ 3);
  assign w80[8] = |(datain[279:276] ^ 13);
  assign w80[9] = |(datain[275:272] ^ 2);
  assign w80[10] = |(datain[271:268] ^ 12);
  assign w80[11] = |(datain[267:264] ^ 13);
  assign w80[12] = |(datain[263:260] ^ 2);
  assign w80[13] = |(datain[259:256] ^ 1);
  assign w80[14] = |(datain[255:252] ^ 11);
  assign w80[15] = |(datain[251:248] ^ 4);
  assign w80[16] = |(datain[247:244] ^ 4);
  assign w80[17] = |(datain[243:240] ^ 0);
  assign w80[18] = |(datain[239:236] ^ 11);
  assign w80[19] = |(datain[235:232] ^ 9);
  assign w80[20] = |(datain[231:228] ^ 0);
  assign w80[21] = |(datain[227:224] ^ 3);
  assign w80[22] = |(datain[223:220] ^ 0);
  assign w80[23] = |(datain[219:216] ^ 0);
  assign w80[24] = |(datain[215:212] ^ 11);
  assign w80[25] = |(datain[211:208] ^ 10);
  assign w80[26] = |(datain[207:204] ^ 2);
  assign w80[27] = |(datain[203:200] ^ 12);
  assign w80[28] = |(datain[199:196] ^ 15);
  assign w80[29] = |(datain[195:192] ^ 11);
  assign w80[30] = |(datain[191:188] ^ 12);
  assign w80[31] = |(datain[187:184] ^ 13);
  assign w80[32] = |(datain[183:180] ^ 2);
  assign w80[33] = |(datain[179:176] ^ 1);
  assign w80[34] = |(datain[175:172] ^ 11);
  assign w80[35] = |(datain[171:168] ^ 8);
  assign w80[36] = |(datain[167:164] ^ 0);
  assign w80[37] = |(datain[163:160] ^ 1);
  assign w80[38] = |(datain[159:156] ^ 5);
  assign w80[39] = |(datain[155:152] ^ 7);
  assign w80[40] = |(datain[151:148] ^ 2);
  assign w80[41] = |(datain[147:144] ^ 14);
  assign w80[42] = |(datain[143:140] ^ 8);
  assign w80[43] = |(datain[139:136] ^ 11);
  assign w80[44] = |(datain[135:132] ^ 1);
  assign w80[45] = |(datain[131:128] ^ 6);
  assign w80[46] = |(datain[127:124] ^ 12);
  assign w80[47] = |(datain[123:120] ^ 10);
  assign w80[48] = |(datain[119:116] ^ 15);
  assign w80[49] = |(datain[115:112] ^ 10);
  assign w80[50] = |(datain[111:108] ^ 2);
  assign w80[51] = |(datain[107:104] ^ 14);
  assign w80[52] = |(datain[103:100] ^ 8);
  assign w80[53] = |(datain[99:96] ^ 11);
  assign w80[54] = |(datain[95:92] ^ 0);
  assign w80[55] = |(datain[91:88] ^ 14);
  assign w80[56] = |(datain[87:84] ^ 12);
  assign w80[57] = |(datain[83:80] ^ 8);
  assign w80[58] = |(datain[79:76] ^ 15);
  assign w80[59] = |(datain[75:72] ^ 10);
  assign w80[60] = |(datain[71:68] ^ 8);
  assign w80[61] = |(datain[67:64] ^ 0);
  assign w80[62] = |(datain[63:60] ^ 14);
  assign w80[63] = |(datain[59:56] ^ 1);
  assign w80[64] = |(datain[55:52] ^ 14);
  assign w80[65] = |(datain[51:48] ^ 0);
  assign w80[66] = |(datain[47:44] ^ 8);
  assign w80[67] = |(datain[43:40] ^ 0);
  assign w80[68] = |(datain[39:36] ^ 12);
  assign w80[69] = |(datain[35:32] ^ 9);
  assign w80[70] = |(datain[31:28] ^ 0);
  assign w80[71] = |(datain[27:24] ^ 3);
  assign w80[72] = |(datain[23:20] ^ 12);
  assign w80[73] = |(datain[19:16] ^ 13);
  assign comp[80] = ~(|w80);
  wire [74-1:0] w81;
  assign w81[0] = |(datain[311:308] ^ 11);
  assign w81[1] = |(datain[307:304] ^ 8);
  assign w81[2] = |(datain[303:300] ^ 0);
  assign w81[3] = |(datain[299:296] ^ 2);
  assign w81[4] = |(datain[295:292] ^ 4);
  assign w81[5] = |(datain[291:288] ^ 2);
  assign w81[6] = |(datain[287:284] ^ 14);
  assign w81[7] = |(datain[283:280] ^ 8);
  assign w81[8] = |(datain[279:276] ^ 4);
  assign w81[9] = |(datain[275:272] ^ 14);
  assign w81[10] = |(datain[271:268] ^ 0);
  assign w81[11] = |(datain[267:264] ^ 0);
  assign w81[12] = |(datain[263:260] ^ 11);
  assign w81[13] = |(datain[259:256] ^ 4);
  assign w81[14] = |(datain[255:252] ^ 4);
  assign w81[15] = |(datain[251:248] ^ 0);
  assign w81[16] = |(datain[247:244] ^ 11);
  assign w81[17] = |(datain[243:240] ^ 10);
  assign w81[18] = |(datain[239:236] ^ 3);
  assign w81[19] = |(datain[235:232] ^ 14);
  assign w81[20] = |(datain[231:228] ^ 15);
  assign w81[21] = |(datain[227:224] ^ 14);
  assign w81[22] = |(datain[223:220] ^ 11);
  assign w81[23] = |(datain[219:216] ^ 9);
  assign w81[24] = |(datain[215:212] ^ 14);
  assign w81[25] = |(datain[211:208] ^ 3);
  assign w81[26] = |(datain[207:204] ^ 0);
  assign w81[27] = |(datain[203:200] ^ 0);
  assign w81[28] = |(datain[199:196] ^ 9);
  assign w81[29] = |(datain[195:192] ^ 0);
  assign w81[30] = |(datain[191:188] ^ 12);
  assign w81[31] = |(datain[187:184] ^ 13);
  assign w81[32] = |(datain[183:180] ^ 2);
  assign w81[33] = |(datain[179:176] ^ 1);
  assign w81[34] = |(datain[175:172] ^ 7);
  assign w81[35] = |(datain[171:168] ^ 2);
  assign w81[36] = |(datain[167:164] ^ 1);
  assign w81[37] = |(datain[163:160] ^ 3);
  assign w81[38] = |(datain[159:156] ^ 11);
  assign w81[39] = |(datain[155:152] ^ 8);
  assign w81[40] = |(datain[151:148] ^ 0);
  assign w81[41] = |(datain[147:144] ^ 0);
  assign w81[42] = |(datain[143:140] ^ 4);
  assign w81[43] = |(datain[139:136] ^ 2);
  assign w81[44] = |(datain[135:132] ^ 14);
  assign w81[45] = |(datain[131:128] ^ 8);
  assign w81[46] = |(datain[127:124] ^ 3);
  assign w81[47] = |(datain[123:120] ^ 11);
  assign w81[48] = |(datain[119:116] ^ 0);
  assign w81[49] = |(datain[115:112] ^ 0);
  assign w81[50] = |(datain[111:108] ^ 11);
  assign w81[51] = |(datain[107:104] ^ 4);
  assign w81[52] = |(datain[103:100] ^ 4);
  assign w81[53] = |(datain[99:96] ^ 0);
  assign w81[54] = |(datain[95:92] ^ 11);
  assign w81[55] = |(datain[91:88] ^ 10);
  assign w81[56] = |(datain[87:84] ^ 0);
  assign w81[57] = |(datain[83:80] ^ 0);
  assign w81[58] = |(datain[79:76] ^ 0);
  assign w81[59] = |(datain[75:72] ^ 1);
  assign w81[60] = |(datain[71:68] ^ 11);
  assign w81[61] = |(datain[67:64] ^ 9);
  assign w81[62] = |(datain[63:60] ^ 14);
  assign w81[63] = |(datain[59:56] ^ 3);
  assign w81[64] = |(datain[55:52] ^ 0);
  assign w81[65] = |(datain[51:48] ^ 0);
  assign w81[66] = |(datain[47:44] ^ 9);
  assign w81[67] = |(datain[43:40] ^ 0);
  assign w81[68] = |(datain[39:36] ^ 12);
  assign w81[69] = |(datain[35:32] ^ 13);
  assign w81[70] = |(datain[31:28] ^ 2);
  assign w81[71] = |(datain[27:24] ^ 1);
  assign w81[72] = |(datain[23:20] ^ 7);
  assign w81[73] = |(datain[19:16] ^ 2);
  assign comp[81] = ~(|w81);
  wire [76-1:0] w82;
  assign w82[0] = |(datain[311:308] ^ 1);
  assign w82[1] = |(datain[307:304] ^ 3);
  assign w82[2] = |(datain[303:300] ^ 11);
  assign w82[3] = |(datain[299:296] ^ 8);
  assign w82[4] = |(datain[295:292] ^ 0);
  assign w82[5] = |(datain[291:288] ^ 0);
  assign w82[6] = |(datain[287:284] ^ 4);
  assign w82[7] = |(datain[283:280] ^ 2);
  assign w82[8] = |(datain[279:276] ^ 14);
  assign w82[9] = |(datain[275:272] ^ 8);
  assign w82[10] = |(datain[271:268] ^ 3);
  assign w82[11] = |(datain[267:264] ^ 11);
  assign w82[12] = |(datain[263:260] ^ 0);
  assign w82[13] = |(datain[259:256] ^ 0);
  assign w82[14] = |(datain[255:252] ^ 11);
  assign w82[15] = |(datain[251:248] ^ 4);
  assign w82[16] = |(datain[247:244] ^ 4);
  assign w82[17] = |(datain[243:240] ^ 0);
  assign w82[18] = |(datain[239:236] ^ 11);
  assign w82[19] = |(datain[235:232] ^ 10);
  assign w82[20] = |(datain[231:228] ^ 0);
  assign w82[21] = |(datain[227:224] ^ 0);
  assign w82[22] = |(datain[223:220] ^ 0);
  assign w82[23] = |(datain[219:216] ^ 1);
  assign w82[24] = |(datain[215:212] ^ 11);
  assign w82[25] = |(datain[211:208] ^ 9);
  assign w82[26] = |(datain[207:204] ^ 14);
  assign w82[27] = |(datain[203:200] ^ 3);
  assign w82[28] = |(datain[199:196] ^ 0);
  assign w82[29] = |(datain[195:192] ^ 0);
  assign w82[30] = |(datain[191:188] ^ 9);
  assign w82[31] = |(datain[187:184] ^ 0);
  assign w82[32] = |(datain[183:180] ^ 12);
  assign w82[33] = |(datain[179:176] ^ 13);
  assign w82[34] = |(datain[175:172] ^ 2);
  assign w82[35] = |(datain[171:168] ^ 1);
  assign w82[36] = |(datain[167:164] ^ 7);
  assign w82[37] = |(datain[163:160] ^ 2);
  assign w82[38] = |(datain[159:156] ^ 0);
  assign w82[39] = |(datain[155:152] ^ 0);
  assign w82[40] = |(datain[151:148] ^ 11);
  assign w82[41] = |(datain[147:144] ^ 4);
  assign w82[42] = |(datain[143:140] ^ 3);
  assign w82[43] = |(datain[139:136] ^ 14);
  assign w82[44] = |(datain[135:132] ^ 12);
  assign w82[45] = |(datain[131:128] ^ 13);
  assign w82[46] = |(datain[127:124] ^ 2);
  assign w82[47] = |(datain[123:120] ^ 1);
  assign w82[48] = |(datain[119:116] ^ 11);
  assign w82[49] = |(datain[115:112] ^ 14);
  assign w82[50] = |(datain[111:108] ^ 10);
  assign w82[51] = |(datain[107:104] ^ 12);
  assign w82[52] = |(datain[103:100] ^ 0);
  assign w82[53] = |(datain[99:96] ^ 1);
  assign w82[54] = |(datain[95:92] ^ 11);
  assign w82[55] = |(datain[91:88] ^ 15);
  assign w82[56] = |(datain[87:84] ^ 3);
  assign w82[57] = |(datain[83:80] ^ 14);
  assign w82[58] = |(datain[79:76] ^ 15);
  assign w82[59] = |(datain[75:72] ^ 15);
  assign w82[60] = |(datain[71:68] ^ 5);
  assign w82[61] = |(datain[67:64] ^ 7);
  assign w82[62] = |(datain[63:60] ^ 11);
  assign w82[63] = |(datain[59:56] ^ 9);
  assign w82[64] = |(datain[55:52] ^ 1);
  assign w82[65] = |(datain[51:48] ^ 9);
  assign w82[66] = |(datain[47:44] ^ 0);
  assign w82[67] = |(datain[43:40] ^ 0);
  assign w82[68] = |(datain[39:36] ^ 9);
  assign w82[69] = |(datain[35:32] ^ 0);
  assign w82[70] = |(datain[31:28] ^ 15);
  assign w82[71] = |(datain[27:24] ^ 12);
  assign w82[72] = |(datain[23:20] ^ 15);
  assign w82[73] = |(datain[19:16] ^ 3);
  assign w82[74] = |(datain[15:12] ^ 10);
  assign w82[75] = |(datain[11:8] ^ 4);
  assign comp[82] = ~(|w82);
  wire [76-1:0] w83;
  assign w83[0] = |(datain[311:308] ^ 8);
  assign w83[1] = |(datain[307:304] ^ 3);
  assign w83[2] = |(datain[303:300] ^ 12);
  assign w83[3] = |(datain[299:296] ^ 0);
  assign w83[4] = |(datain[295:292] ^ 0);
  assign w83[5] = |(datain[291:288] ^ 9);
  assign w83[6] = |(datain[287:284] ^ 8);
  assign w83[7] = |(datain[283:280] ^ 9);
  assign w83[8] = |(datain[279:276] ^ 8);
  assign w83[9] = |(datain[275:272] ^ 6);
  assign w83[10] = |(datain[271:268] ^ 0);
  assign w83[11] = |(datain[267:264] ^ 10);
  assign w83[12] = |(datain[263:260] ^ 0);
  assign w83[13] = |(datain[259:256] ^ 1);
  assign w83[14] = |(datain[255:252] ^ 8);
  assign w83[15] = |(datain[251:248] ^ 13);
  assign w83[16] = |(datain[247:244] ^ 9);
  assign w83[17] = |(datain[243:240] ^ 6);
  assign w83[18] = |(datain[239:236] ^ 0);
  assign w83[19] = |(datain[235:232] ^ 9);
  assign w83[20] = |(datain[231:228] ^ 0);
  assign w83[21] = |(datain[227:224] ^ 1);
  assign w83[22] = |(datain[223:220] ^ 11);
  assign w83[23] = |(datain[219:216] ^ 4);
  assign w83[24] = |(datain[215:212] ^ 4);
  assign w83[25] = |(datain[211:208] ^ 0);
  assign w83[26] = |(datain[207:204] ^ 11);
  assign w83[27] = |(datain[203:200] ^ 9);
  assign w83[28] = |(datain[199:196] ^ 0);
  assign w83[29] = |(datain[195:192] ^ 3);
  assign w83[30] = |(datain[191:188] ^ 0);
  assign w83[31] = |(datain[187:184] ^ 0);
  assign w83[32] = |(datain[183:180] ^ 12);
  assign w83[33] = |(datain[179:176] ^ 13);
  assign w83[34] = |(datain[175:172] ^ 2);
  assign w83[35] = |(datain[171:168] ^ 1);
  assign w83[36] = |(datain[167:164] ^ 11);
  assign w83[37] = |(datain[163:160] ^ 8);
  assign w83[38] = |(datain[159:156] ^ 0);
  assign w83[39] = |(datain[155:152] ^ 2);
  assign w83[40] = |(datain[151:148] ^ 4);
  assign w83[41] = |(datain[147:144] ^ 2);
  assign w83[42] = |(datain[143:140] ^ 14);
  assign w83[43] = |(datain[139:136] ^ 8);
  assign w83[44] = |(datain[135:132] ^ 2);
  assign w83[45] = |(datain[131:128] ^ 6);
  assign w83[46] = |(datain[127:124] ^ 0);
  assign w83[47] = |(datain[123:120] ^ 0);
  assign w83[48] = |(datain[119:116] ^ 8);
  assign w83[49] = |(datain[115:112] ^ 13);
  assign w83[50] = |(datain[111:108] ^ 9);
  assign w83[51] = |(datain[107:104] ^ 6);
  assign w83[52] = |(datain[103:100] ^ 0);
  assign w83[53] = |(datain[99:96] ^ 3);
  assign w83[54] = |(datain[95:92] ^ 0);
  assign w83[55] = |(datain[91:88] ^ 1);
  assign w83[56] = |(datain[87:84] ^ 11);
  assign w83[57] = |(datain[83:80] ^ 4);
  assign w83[58] = |(datain[79:76] ^ 4);
  assign w83[59] = |(datain[75:72] ^ 0);
  assign w83[60] = |(datain[71:68] ^ 11);
  assign w83[61] = |(datain[67:64] ^ 9);
  assign w83[62] = |(datain[63:60] ^ 11);
  assign w83[63] = |(datain[59:56] ^ 2);
  assign w83[64] = |(datain[55:52] ^ 0);
  assign w83[65] = |(datain[51:48] ^ 0);
  assign w83[66] = |(datain[47:44] ^ 12);
  assign w83[67] = |(datain[43:40] ^ 13);
  assign w83[68] = |(datain[39:36] ^ 2);
  assign w83[69] = |(datain[35:32] ^ 1);
  assign w83[70] = |(datain[31:28] ^ 11);
  assign w83[71] = |(datain[27:24] ^ 8);
  assign w83[72] = |(datain[23:20] ^ 0);
  assign w83[73] = |(datain[19:16] ^ 1);
  assign w83[74] = |(datain[15:12] ^ 5);
  assign w83[75] = |(datain[11:8] ^ 7);
  assign comp[83] = ~(|w83);
  wire [76-1:0] w84;
  assign w84[0] = |(datain[311:308] ^ 12);
  assign w84[1] = |(datain[307:304] ^ 9);
  assign w84[2] = |(datain[303:300] ^ 14);
  assign w84[3] = |(datain[299:296] ^ 8);
  assign w84[4] = |(datain[295:292] ^ 0);
  assign w84[5] = |(datain[291:288] ^ 8);
  assign w84[6] = |(datain[287:284] ^ 0);
  assign w84[7] = |(datain[283:280] ^ 0);
  assign w84[8] = |(datain[279:276] ^ 8);
  assign w84[9] = |(datain[275:272] ^ 11);
  assign w84[10] = |(datain[271:268] ^ 13);
  assign w84[11] = |(datain[267:264] ^ 0);
  assign w84[12] = |(datain[263:260] ^ 11);
  assign w84[13] = |(datain[259:256] ^ 4);
  assign w84[14] = |(datain[255:252] ^ 4);
  assign w84[15] = |(datain[251:248] ^ 0);
  assign w84[16] = |(datain[247:244] ^ 11);
  assign w84[17] = |(datain[243:240] ^ 9);
  assign w84[18] = |(datain[239:236] ^ 0);
  assign w84[19] = |(datain[235:232] ^ 3);
  assign w84[20] = |(datain[231:228] ^ 0);
  assign w84[21] = |(datain[227:224] ^ 0);
  assign w84[22] = |(datain[223:220] ^ 12);
  assign w84[23] = |(datain[219:216] ^ 3);
  assign w84[24] = |(datain[215:212] ^ 9);
  assign w84[25] = |(datain[211:208] ^ 12);
  assign w84[26] = |(datain[207:204] ^ 2);
  assign w84[27] = |(datain[203:200] ^ 14);
  assign w84[28] = |(datain[199:196] ^ 15);
  assign w84[29] = |(datain[195:192] ^ 15);
  assign w84[30] = |(datain[191:188] ^ 9);
  assign w84[31] = |(datain[187:184] ^ 14);
  assign w84[32] = |(datain[183:180] ^ 8);
  assign w84[33] = |(datain[179:176] ^ 7);
  assign w84[34] = |(datain[175:172] ^ 0);
  assign w84[35] = |(datain[171:168] ^ 2);
  assign w84[36] = |(datain[167:164] ^ 12);
  assign w84[37] = |(datain[163:160] ^ 3);
  assign w84[38] = |(datain[159:156] ^ 3);
  assign w84[39] = |(datain[155:152] ^ 3);
  assign w84[40] = |(datain[151:148] ^ 12);
  assign w84[41] = |(datain[147:144] ^ 0);
  assign w84[42] = |(datain[143:140] ^ 8);
  assign w84[43] = |(datain[139:136] ^ 14);
  assign w84[44] = |(datain[135:132] ^ 13);
  assign w84[45] = |(datain[131:128] ^ 8);
  assign w84[46] = |(datain[127:124] ^ 8);
  assign w84[47] = |(datain[123:120] ^ 11);
  assign w84[48] = |(datain[119:116] ^ 3);
  assign w84[49] = |(datain[115:112] ^ 6);
  assign w84[50] = |(datain[111:108] ^ 0);
  assign w84[51] = |(datain[107:104] ^ 4);
  assign w84[52] = |(datain[103:100] ^ 0);
  assign w84[53] = |(datain[99:96] ^ 0);
  assign w84[54] = |(datain[95:92] ^ 8);
  assign w84[55] = |(datain[91:88] ^ 11);
  assign w84[56] = |(datain[87:84] ^ 1);
  assign w84[57] = |(datain[83:80] ^ 14);
  assign w84[58] = |(datain[79:76] ^ 0);
  assign w84[59] = |(datain[75:72] ^ 6);
  assign w84[60] = |(datain[71:68] ^ 0);
  assign w84[61] = |(datain[67:64] ^ 0);
  assign w84[62] = |(datain[63:60] ^ 8);
  assign w84[63] = |(datain[59:56] ^ 14);
  assign w84[64] = |(datain[55:52] ^ 12);
  assign w84[65] = |(datain[51:48] ^ 3);
  assign w84[66] = |(datain[47:44] ^ 5);
  assign w84[67] = |(datain[43:40] ^ 0);
  assign w84[68] = |(datain[39:36] ^ 9);
  assign w84[69] = |(datain[35:32] ^ 13);
  assign w84[70] = |(datain[31:28] ^ 10);
  assign w84[71] = |(datain[27:24] ^ 1);
  assign w84[72] = |(datain[23:20] ^ 10);
  assign w84[73] = |(datain[19:16] ^ 14);
  assign w84[74] = |(datain[15:12] ^ 0);
  assign w84[75] = |(datain[11:8] ^ 0);
  assign comp[84] = ~(|w84);
  wire [76-1:0] w85;
  assign w85[0] = |(datain[311:308] ^ 3);
  assign w85[1] = |(datain[307:304] ^ 5);
  assign w85[2] = |(datain[303:300] ^ 10);
  assign w85[3] = |(datain[299:296] ^ 13);
  assign w85[4] = |(datain[295:292] ^ 0);
  assign w85[5] = |(datain[291:288] ^ 0);
  assign w85[6] = |(datain[287:284] ^ 8);
  assign w85[7] = |(datain[283:280] ^ 9);
  assign w85[8] = |(datain[279:276] ^ 0);
  assign w85[9] = |(datain[275:272] ^ 5);
  assign w85[10] = |(datain[271:268] ^ 4);
  assign w85[11] = |(datain[267:264] ^ 7);
  assign w85[12] = |(datain[263:260] ^ 4);
  assign w85[13] = |(datain[259:256] ^ 7);
  assign w85[14] = |(datain[255:252] ^ 14);
  assign w85[15] = |(datain[251:248] ^ 2);
  assign w85[16] = |(datain[247:244] ^ 15);
  assign w85[17] = |(datain[243:240] ^ 0);
  assign w85[18] = |(datain[239:236] ^ 14);
  assign w85[19] = |(datain[235:232] ^ 8);
  assign w85[20] = |(datain[231:228] ^ 3);
  assign w85[21] = |(datain[227:224] ^ 7);
  assign w85[22] = |(datain[223:220] ^ 0);
  assign w85[23] = |(datain[219:216] ^ 0);
  assign w85[24] = |(datain[215:212] ^ 11);
  assign w85[25] = |(datain[211:208] ^ 4);
  assign w85[26] = |(datain[207:204] ^ 4);
  assign w85[27] = |(datain[203:200] ^ 0);
  assign w85[28] = |(datain[199:196] ^ 5);
  assign w85[29] = |(datain[195:192] ^ 10);
  assign w85[30] = |(datain[191:188] ^ 5);
  assign w85[31] = |(datain[187:184] ^ 9);
  assign w85[32] = |(datain[183:180] ^ 12);
  assign w85[33] = |(datain[179:176] ^ 13);
  assign w85[34] = |(datain[175:172] ^ 2);
  assign w85[35] = |(datain[171:168] ^ 1);
  assign w85[36] = |(datain[167:164] ^ 14);
  assign w85[37] = |(datain[163:160] ^ 8);
  assign w85[38] = |(datain[159:156] ^ 3);
  assign w85[39] = |(datain[155:152] ^ 8);
  assign w85[40] = |(datain[151:148] ^ 0);
  assign w85[41] = |(datain[147:144] ^ 0);
  assign w85[42] = |(datain[143:140] ^ 11);
  assign w85[43] = |(datain[139:136] ^ 4);
  assign w85[44] = |(datain[135:132] ^ 4);
  assign w85[45] = |(datain[131:128] ^ 0);
  assign w85[46] = |(datain[127:124] ^ 11);
  assign w85[47] = |(datain[123:120] ^ 9);
  assign w85[48] = |(datain[119:116] ^ 4);
  assign w85[49] = |(datain[115:112] ^ 4);
  assign w85[50] = |(datain[111:108] ^ 0);
  assign w85[51] = |(datain[107:104] ^ 2);
  assign w85[52] = |(datain[103:100] ^ 9);
  assign w85[53] = |(datain[99:96] ^ 0);
  assign w85[54] = |(datain[95:92] ^ 11);
  assign w85[55] = |(datain[91:88] ^ 10);
  assign w85[56] = |(datain[87:84] ^ 0);
  assign w85[57] = |(datain[83:80] ^ 0);
  assign w85[58] = |(datain[79:76] ^ 0);
  assign w85[59] = |(datain[75:72] ^ 1);
  assign w85[60] = |(datain[71:68] ^ 12);
  assign w85[61] = |(datain[67:64] ^ 13);
  assign w85[62] = |(datain[63:60] ^ 2);
  assign w85[63] = |(datain[59:56] ^ 1);
  assign w85[64] = |(datain[55:52] ^ 11);
  assign w85[65] = |(datain[51:48] ^ 8);
  assign w85[66] = |(datain[47:44] ^ 0);
  assign w85[67] = |(datain[43:40] ^ 1);
  assign w85[68] = |(datain[39:36] ^ 5);
  assign w85[69] = |(datain[35:32] ^ 7);
  assign w85[70] = |(datain[31:28] ^ 8);
  assign w85[71] = |(datain[27:24] ^ 11);
  assign w85[72] = |(datain[23:20] ^ 3);
  assign w85[73] = |(datain[19:16] ^ 6);
  assign w85[74] = |(datain[15:12] ^ 15);
  assign w85[75] = |(datain[11:8] ^ 13);
  assign comp[85] = ~(|w85);
  wire [74-1:0] w86;
  assign w86[0] = |(datain[311:308] ^ 13);
  assign w86[1] = |(datain[307:304] ^ 2);
  assign w86[2] = |(datain[303:300] ^ 11);
  assign w86[3] = |(datain[299:296] ^ 8);
  assign w86[4] = |(datain[295:292] ^ 0);
  assign w86[5] = |(datain[291:288] ^ 0);
  assign w86[6] = |(datain[287:284] ^ 4);
  assign w86[7] = |(datain[283:280] ^ 2);
  assign w86[8] = |(datain[279:276] ^ 12);
  assign w86[9] = |(datain[275:272] ^ 13);
  assign w86[10] = |(datain[271:268] ^ 2);
  assign w86[11] = |(datain[267:264] ^ 1);
  assign w86[12] = |(datain[263:260] ^ 11);
  assign w86[13] = |(datain[259:256] ^ 9);
  assign w86[14] = |(datain[255:252] ^ 2);
  assign w86[15] = |(datain[251:248] ^ 0);
  assign w86[16] = |(datain[247:244] ^ 0);
  assign w86[17] = |(datain[243:240] ^ 0);
  assign w86[18] = |(datain[239:236] ^ 8);
  assign w86[19] = |(datain[235:232] ^ 13);
  assign w86[20] = |(datain[231:228] ^ 9);
  assign w86[21] = |(datain[227:224] ^ 6);
  assign w86[22] = |(datain[223:220] ^ 13);
  assign w86[23] = |(datain[219:216] ^ 11);
  assign w86[24] = |(datain[215:212] ^ 0);
  assign w86[25] = |(datain[211:208] ^ 3);
  assign w86[26] = |(datain[207:204] ^ 11);
  assign w86[27] = |(datain[203:200] ^ 4);
  assign w86[28] = |(datain[199:196] ^ 4);
  assign w86[29] = |(datain[195:192] ^ 0);
  assign w86[30] = |(datain[191:188] ^ 12);
  assign w86[31] = |(datain[187:184] ^ 13);
  assign w86[32] = |(datain[183:180] ^ 2);
  assign w86[33] = |(datain[179:176] ^ 1);
  assign w86[34] = |(datain[175:172] ^ 7);
  assign w86[35] = |(datain[171:168] ^ 2);
  assign w86[36] = |(datain[167:164] ^ 0);
  assign w86[37] = |(datain[163:160] ^ 13);
  assign w86[38] = |(datain[159:156] ^ 8);
  assign w86[39] = |(datain[155:152] ^ 11);
  assign w86[40] = |(datain[151:148] ^ 8);
  assign w86[41] = |(datain[147:144] ^ 14);
  assign w86[42] = |(datain[143:140] ^ 1);
  assign w86[43] = |(datain[139:136] ^ 3);
  assign w86[44] = |(datain[135:132] ^ 0);
  assign w86[45] = |(datain[131:128] ^ 4);
  assign w86[46] = |(datain[127:124] ^ 8);
  assign w86[47] = |(datain[123:120] ^ 11);
  assign w86[48] = |(datain[119:116] ^ 9);
  assign w86[49] = |(datain[115:112] ^ 6);
  assign w86[50] = |(datain[111:108] ^ 1);
  assign w86[51] = |(datain[107:104] ^ 5);
  assign w86[52] = |(datain[103:100] ^ 0);
  assign w86[53] = |(datain[99:96] ^ 4);
  assign w86[54] = |(datain[95:92] ^ 11);
  assign w86[55] = |(datain[91:88] ^ 8);
  assign w86[56] = |(datain[87:84] ^ 0);
  assign w86[57] = |(datain[83:80] ^ 1);
  assign w86[58] = |(datain[79:76] ^ 5);
  assign w86[59] = |(datain[75:72] ^ 7);
  assign w86[60] = |(datain[71:68] ^ 12);
  assign w86[61] = |(datain[67:64] ^ 13);
  assign w86[62] = |(datain[63:60] ^ 2);
  assign w86[63] = |(datain[59:56] ^ 1);
  assign w86[64] = |(datain[55:52] ^ 11);
  assign w86[65] = |(datain[51:48] ^ 4);
  assign w86[66] = |(datain[47:44] ^ 3);
  assign w86[67] = |(datain[43:40] ^ 14);
  assign w86[68] = |(datain[39:36] ^ 12);
  assign w86[69] = |(datain[35:32] ^ 13);
  assign w86[70] = |(datain[31:28] ^ 2);
  assign w86[71] = |(datain[27:24] ^ 1);
  assign w86[72] = |(datain[23:20] ^ 8);
  assign w86[73] = |(datain[19:16] ^ 13);
  assign comp[86] = ~(|w86);
  wire [74-1:0] w87;
  assign w87[0] = |(datain[311:308] ^ 13);
  assign w87[1] = |(datain[307:304] ^ 2);
  assign w87[2] = |(datain[303:300] ^ 11);
  assign w87[3] = |(datain[299:296] ^ 8);
  assign w87[4] = |(datain[295:292] ^ 0);
  assign w87[5] = |(datain[291:288] ^ 2);
  assign w87[6] = |(datain[287:284] ^ 4);
  assign w87[7] = |(datain[283:280] ^ 2);
  assign w87[8] = |(datain[279:276] ^ 12);
  assign w87[9] = |(datain[275:272] ^ 13);
  assign w87[10] = |(datain[271:268] ^ 2);
  assign w87[11] = |(datain[267:264] ^ 1);
  assign w87[12] = |(datain[263:260] ^ 11);
  assign w87[13] = |(datain[259:256] ^ 9);
  assign w87[14] = |(datain[255:252] ^ 1);
  assign w87[15] = |(datain[251:248] ^ 7);
  assign w87[16] = |(datain[247:244] ^ 0);
  assign w87[17] = |(datain[243:240] ^ 0);
  assign w87[18] = |(datain[239:236] ^ 8);
  assign w87[19] = |(datain[235:232] ^ 13);
  assign w87[20] = |(datain[231:228] ^ 9);
  assign w87[21] = |(datain[227:224] ^ 6);
  assign w87[22] = |(datain[223:220] ^ 0);
  assign w87[23] = |(datain[219:216] ^ 0);
  assign w87[24] = |(datain[215:212] ^ 0);
  assign w87[25] = |(datain[211:208] ^ 1);
  assign w87[26] = |(datain[207:204] ^ 11);
  assign w87[27] = |(datain[203:200] ^ 4);
  assign w87[28] = |(datain[199:196] ^ 4);
  assign w87[29] = |(datain[195:192] ^ 0);
  assign w87[30] = |(datain[191:188] ^ 12);
  assign w87[31] = |(datain[187:184] ^ 13);
  assign w87[32] = |(datain[183:180] ^ 2);
  assign w87[33] = |(datain[179:176] ^ 1);
  assign w87[34] = |(datain[175:172] ^ 7);
  assign w87[35] = |(datain[171:168] ^ 2);
  assign w87[36] = |(datain[167:164] ^ 3);
  assign w87[37] = |(datain[163:160] ^ 4);
  assign w87[38] = |(datain[159:156] ^ 1);
  assign w87[39] = |(datain[155:152] ^ 14);
  assign w87[40] = |(datain[151:148] ^ 8);
  assign w87[41] = |(datain[147:144] ^ 12);
  assign w87[42] = |(datain[143:140] ^ 12);
  assign w87[43] = |(datain[139:136] ^ 0);
  assign w87[44] = |(datain[135:132] ^ 8);
  assign w87[45] = |(datain[131:128] ^ 14);
  assign w87[46] = |(datain[127:124] ^ 13);
  assign w87[47] = |(datain[123:120] ^ 8);
  assign w87[48] = |(datain[119:116] ^ 11);
  assign w87[49] = |(datain[115:112] ^ 9);
  assign w87[50] = |(datain[111:108] ^ 12);
  assign w87[51] = |(datain[107:104] ^ 4);
  assign w87[52] = |(datain[103:100] ^ 0);
  assign w87[53] = |(datain[99:96] ^ 2);
  assign w87[54] = |(datain[95:92] ^ 3);
  assign w87[55] = |(datain[91:88] ^ 3);
  assign w87[56] = |(datain[87:84] ^ 13);
  assign w87[57] = |(datain[83:80] ^ 2);
  assign w87[58] = |(datain[79:76] ^ 11);
  assign w87[59] = |(datain[75:72] ^ 4);
  assign w87[60] = |(datain[71:68] ^ 4);
  assign w87[61] = |(datain[67:64] ^ 0);
  assign w87[62] = |(datain[63:60] ^ 12);
  assign w87[63] = |(datain[59:56] ^ 13);
  assign w87[64] = |(datain[55:52] ^ 2);
  assign w87[65] = |(datain[51:48] ^ 1);
  assign w87[66] = |(datain[47:44] ^ 1);
  assign w87[67] = |(datain[43:40] ^ 15);
  assign w87[68] = |(datain[39:36] ^ 7);
  assign w87[69] = |(datain[35:32] ^ 2);
  assign w87[70] = |(datain[31:28] ^ 2);
  assign w87[71] = |(datain[27:24] ^ 3);
  assign w87[72] = |(datain[23:20] ^ 3);
  assign w87[73] = |(datain[19:16] ^ 3);
  assign comp[87] = ~(|w87);
  wire [74-1:0] w88;
  assign w88[0] = |(datain[311:308] ^ 2);
  assign w88[1] = |(datain[307:304] ^ 8);
  assign w88[2] = |(datain[303:300] ^ 10);
  assign w88[3] = |(datain[299:296] ^ 3);
  assign w88[4] = |(datain[295:292] ^ 8);
  assign w88[5] = |(datain[291:288] ^ 4);
  assign w88[6] = |(datain[287:284] ^ 0);
  assign w88[7] = |(datain[283:280] ^ 0);
  assign w88[8] = |(datain[279:276] ^ 11);
  assign w88[9] = |(datain[275:272] ^ 8);
  assign w88[10] = |(datain[271:268] ^ 0);
  assign w88[11] = |(datain[267:264] ^ 0);
  assign w88[12] = |(datain[263:260] ^ 5);
  assign w88[13] = |(datain[259:256] ^ 7);
  assign w88[14] = |(datain[255:252] ^ 12);
  assign w88[15] = |(datain[251:248] ^ 12);
  assign w88[16] = |(datain[247:244] ^ 5);
  assign w88[17] = |(datain[243:240] ^ 1);
  assign w88[18] = |(datain[239:236] ^ 5);
  assign w88[19] = |(datain[235:232] ^ 2);
  assign w88[20] = |(datain[231:228] ^ 11);
  assign w88[21] = |(datain[227:224] ^ 9);
  assign w88[22] = |(datain[223:220] ^ 7);
  assign w88[23] = |(datain[219:216] ^ 2);
  assign w88[24] = |(datain[215:212] ^ 0);
  assign w88[25] = |(datain[211:208] ^ 1);
  assign w88[26] = |(datain[207:204] ^ 11);
  assign w88[27] = |(datain[203:200] ^ 4);
  assign w88[28] = |(datain[199:196] ^ 4);
  assign w88[29] = |(datain[195:192] ^ 0);
  assign w88[30] = |(datain[191:188] ^ 9);
  assign w88[31] = |(datain[187:184] ^ 9);
  assign w88[32] = |(datain[183:180] ^ 12);
  assign w88[33] = |(datain[179:176] ^ 12);
  assign w88[34] = |(datain[175:172] ^ 7);
  assign w88[35] = |(datain[171:168] ^ 2);
  assign w88[36] = |(datain[167:164] ^ 1);
  assign w88[37] = |(datain[163:160] ^ 0);
  assign w88[38] = |(datain[159:156] ^ 11);
  assign w88[39] = |(datain[155:152] ^ 8);
  assign w88[40] = |(datain[151:148] ^ 0);
  assign w88[41] = |(datain[147:144] ^ 0);
  assign w88[42] = |(datain[143:140] ^ 4);
  assign w88[43] = |(datain[139:136] ^ 2);
  assign w88[44] = |(datain[135:132] ^ 3);
  assign w88[45] = |(datain[131:128] ^ 3);
  assign w88[46] = |(datain[127:124] ^ 12);
  assign w88[47] = |(datain[123:120] ^ 9);
  assign w88[48] = |(datain[119:116] ^ 9);
  assign w88[49] = |(datain[115:112] ^ 9);
  assign w88[50] = |(datain[111:108] ^ 12);
  assign w88[51] = |(datain[107:104] ^ 12);
  assign w88[52] = |(datain[103:100] ^ 11);
  assign w88[53] = |(datain[99:96] ^ 9);
  assign w88[54] = |(datain[95:92] ^ 0);
  assign w88[55] = |(datain[91:88] ^ 4);
  assign w88[56] = |(datain[87:84] ^ 0);
  assign w88[57] = |(datain[83:80] ^ 0);
  assign w88[58] = |(datain[79:76] ^ 11);
  assign w88[59] = |(datain[75:72] ^ 10);
  assign w88[60] = |(datain[71:68] ^ 8);
  assign w88[61] = |(datain[67:64] ^ 2);
  assign w88[62] = |(datain[63:60] ^ 0);
  assign w88[63] = |(datain[59:56] ^ 0);
  assign w88[64] = |(datain[55:52] ^ 11);
  assign w88[65] = |(datain[51:48] ^ 4);
  assign w88[66] = |(datain[47:44] ^ 4);
  assign w88[67] = |(datain[43:40] ^ 0);
  assign w88[68] = |(datain[39:36] ^ 12);
  assign w88[69] = |(datain[35:32] ^ 12);
  assign w88[70] = |(datain[31:28] ^ 11);
  assign w88[71] = |(datain[27:24] ^ 8);
  assign w88[72] = |(datain[23:20] ^ 0);
  assign w88[73] = |(datain[19:16] ^ 1);
  assign comp[88] = ~(|w88);
  wire [76-1:0] w89;
  assign w89[0] = |(datain[311:308] ^ 11);
  assign w89[1] = |(datain[307:304] ^ 8);
  assign w89[2] = |(datain[303:300] ^ 0);
  assign w89[3] = |(datain[299:296] ^ 0);
  assign w89[4] = |(datain[295:292] ^ 4);
  assign w89[5] = |(datain[291:288] ^ 2);
  assign w89[6] = |(datain[287:284] ^ 3);
  assign w89[7] = |(datain[283:280] ^ 3);
  assign w89[8] = |(datain[279:276] ^ 12);
  assign w89[9] = |(datain[275:272] ^ 9);
  assign w89[10] = |(datain[271:268] ^ 3);
  assign w89[11] = |(datain[267:264] ^ 3);
  assign w89[12] = |(datain[263:260] ^ 13);
  assign w89[13] = |(datain[259:256] ^ 2);
  assign w89[14] = |(datain[255:252] ^ 12);
  assign w89[15] = |(datain[251:248] ^ 13);
  assign w89[16] = |(datain[247:244] ^ 0);
  assign w89[17] = |(datain[243:240] ^ 1);
  assign w89[18] = |(datain[239:236] ^ 11);
  assign w89[19] = |(datain[235:232] ^ 4);
  assign w89[20] = |(datain[231:228] ^ 4);
  assign w89[21] = |(datain[227:224] ^ 0);
  assign w89[22] = |(datain[223:220] ^ 11);
  assign w89[23] = |(datain[219:216] ^ 10);
  assign w89[24] = |(datain[215:212] ^ 4);
  assign w89[25] = |(datain[211:208] ^ 3);
  assign w89[26] = |(datain[207:204] ^ 0);
  assign w89[27] = |(datain[203:200] ^ 5);
  assign w89[28] = |(datain[199:196] ^ 11);
  assign w89[29] = |(datain[195:192] ^ 9);
  assign w89[30] = |(datain[191:188] ^ 0);
  assign w89[31] = |(datain[187:184] ^ 3);
  assign w89[32] = |(datain[183:180] ^ 0);
  assign w89[33] = |(datain[179:176] ^ 0);
  assign w89[34] = |(datain[175:172] ^ 12);
  assign w89[35] = |(datain[171:168] ^ 12);
  assign w89[36] = |(datain[167:164] ^ 5);
  assign w89[37] = |(datain[163:160] ^ 10);
  assign w89[38] = |(datain[159:156] ^ 5);
  assign w89[39] = |(datain[155:152] ^ 9);
  assign w89[40] = |(datain[151:148] ^ 11);
  assign w89[41] = |(datain[147:144] ^ 8);
  assign w89[42] = |(datain[143:140] ^ 0);
  assign w89[43] = |(datain[139:136] ^ 1);
  assign w89[44] = |(datain[135:132] ^ 5);
  assign w89[45] = |(datain[131:128] ^ 7);
  assign w89[46] = |(datain[127:124] ^ 12);
  assign w89[47] = |(datain[123:120] ^ 13);
  assign w89[48] = |(datain[119:116] ^ 0);
  assign w89[49] = |(datain[115:112] ^ 1);
  assign w89[50] = |(datain[111:108] ^ 11);
  assign w89[51] = |(datain[107:104] ^ 4);
  assign w89[52] = |(datain[103:100] ^ 3);
  assign w89[53] = |(datain[99:96] ^ 14);
  assign w89[54] = |(datain[95:92] ^ 12);
  assign w89[55] = |(datain[91:88] ^ 12);
  assign w89[56] = |(datain[87:84] ^ 11);
  assign w89[57] = |(datain[83:80] ^ 8);
  assign w89[58] = |(datain[79:76] ^ 0);
  assign w89[59] = |(datain[75:72] ^ 1);
  assign w89[60] = |(datain[71:68] ^ 4);
  assign w89[61] = |(datain[67:64] ^ 3);
  assign w89[62] = |(datain[63:60] ^ 5);
  assign w89[63] = |(datain[59:56] ^ 10);
  assign w89[64] = |(datain[55:52] ^ 1);
  assign w89[65] = |(datain[51:48] ^ 15);
  assign w89[66] = |(datain[47:44] ^ 5);
  assign w89[67] = |(datain[43:40] ^ 9);
  assign w89[68] = |(datain[39:36] ^ 12);
  assign w89[69] = |(datain[35:32] ^ 12);
  assign w89[70] = |(datain[31:28] ^ 14);
  assign w89[71] = |(datain[27:24] ^ 9);
  assign w89[72] = |(datain[23:20] ^ 13);
  assign w89[73] = |(datain[19:16] ^ 15);
  assign w89[74] = |(datain[15:12] ^ 15);
  assign w89[75] = |(datain[11:8] ^ 14);
  assign comp[89] = ~(|w89);
  wire [74-1:0] w90;
  assign w90[0] = |(datain[311:308] ^ 15);
  assign w90[1] = |(datain[307:304] ^ 0);
  assign w90[2] = |(datain[303:300] ^ 3);
  assign w90[3] = |(datain[299:296] ^ 13);
  assign w90[4] = |(datain[295:292] ^ 0);
  assign w90[5] = |(datain[291:288] ^ 0);
  assign w90[6] = |(datain[287:284] ^ 15);
  assign w90[7] = |(datain[283:280] ^ 0);
  assign w90[8] = |(datain[279:276] ^ 7);
  assign w90[9] = |(datain[275:272] ^ 5);
  assign w90[10] = |(datain[271:268] ^ 0);
  assign w90[11] = |(datain[267:264] ^ 2);
  assign w90[12] = |(datain[263:260] ^ 14);
  assign w90[13] = |(datain[259:256] ^ 11);
  assign w90[14] = |(datain[255:252] ^ 3);
  assign w90[15] = |(datain[251:248] ^ 3);
  assign w90[16] = |(datain[247:244] ^ 8);
  assign w90[17] = |(datain[243:240] ^ 11);
  assign w90[18] = |(datain[239:236] ^ 13);
  assign w90[19] = |(datain[235:232] ^ 5);
  assign w90[20] = |(datain[231:228] ^ 11);
  assign w90[21] = |(datain[227:224] ^ 9);
  assign w90[22] = |(datain[223:220] ^ 7);
  assign w90[23] = |(datain[219:216] ^ 0);
  assign w90[24] = |(datain[215:212] ^ 0);
  assign w90[25] = |(datain[211:208] ^ 2);
  assign w90[26] = |(datain[207:204] ^ 11);
  assign w90[27] = |(datain[203:200] ^ 4);
  assign w90[28] = |(datain[199:196] ^ 4);
  assign w90[29] = |(datain[195:192] ^ 0);
  assign w90[30] = |(datain[191:188] ^ 12);
  assign w90[31] = |(datain[187:184] ^ 13);
  assign w90[32] = |(datain[183:180] ^ 2);
  assign w90[33] = |(datain[179:176] ^ 1);
  assign w90[34] = |(datain[175:172] ^ 11);
  assign w90[35] = |(datain[171:168] ^ 8);
  assign w90[36] = |(datain[167:164] ^ 0);
  assign w90[37] = |(datain[163:160] ^ 0);
  assign w90[38] = |(datain[159:156] ^ 4);
  assign w90[39] = |(datain[155:152] ^ 2);
  assign w90[40] = |(datain[151:148] ^ 3);
  assign w90[41] = |(datain[147:144] ^ 3);
  assign w90[42] = |(datain[143:140] ^ 12);
  assign w90[43] = |(datain[139:136] ^ 9);
  assign w90[44] = |(datain[135:132] ^ 3);
  assign w90[45] = |(datain[131:128] ^ 3);
  assign w90[46] = |(datain[127:124] ^ 13);
  assign w90[47] = |(datain[123:120] ^ 2);
  assign w90[48] = |(datain[119:116] ^ 12);
  assign w90[49] = |(datain[115:112] ^ 13);
  assign w90[50] = |(datain[111:108] ^ 2);
  assign w90[51] = |(datain[107:104] ^ 1);
  assign w90[52] = |(datain[103:100] ^ 8);
  assign w90[53] = |(datain[99:96] ^ 1);
  assign w90[54] = |(datain[95:92] ^ 12);
  assign w90[55] = |(datain[91:88] ^ 7);
  assign w90[56] = |(datain[87:84] ^ 7);
  assign w90[57] = |(datain[83:80] ^ 0);
  assign w90[58] = |(datain[79:76] ^ 0);
  assign w90[59] = |(datain[75:72] ^ 2);
  assign w90[60] = |(datain[71:68] ^ 12);
  assign w90[61] = |(datain[67:64] ^ 6);
  assign w90[62] = |(datain[63:60] ^ 0);
  assign w90[63] = |(datain[59:56] ^ 5);
  assign w90[64] = |(datain[55:52] ^ 0);
  assign w90[65] = |(datain[51:48] ^ 3);
  assign w90[66] = |(datain[47:44] ^ 12);
  assign w90[67] = |(datain[43:40] ^ 6);
  assign w90[68] = |(datain[39:36] ^ 4);
  assign w90[69] = |(datain[35:32] ^ 5);
  assign w90[70] = |(datain[31:28] ^ 0);
  assign w90[71] = |(datain[27:24] ^ 1);
  assign w90[72] = |(datain[23:20] ^ 0);
  assign w90[73] = |(datain[19:16] ^ 1);
  assign comp[90] = ~(|w90);
  wire [74-1:0] w91;
  assign w91[0] = |(datain[311:308] ^ 8);
  assign w91[1] = |(datain[307:304] ^ 1);
  assign w91[2] = |(datain[303:300] ^ 12);
  assign w91[3] = |(datain[299:296] ^ 5);
  assign w91[4] = |(datain[295:292] ^ 1);
  assign w91[5] = |(datain[291:288] ^ 2);
  assign w91[6] = |(datain[287:284] ^ 0);
  assign w91[7] = |(datain[283:280] ^ 3);
  assign w91[8] = |(datain[279:276] ^ 14);
  assign w91[9] = |(datain[275:272] ^ 8);
  assign w91[10] = |(datain[271:268] ^ 8);
  assign w91[11] = |(datain[267:264] ^ 8);
  assign w91[12] = |(datain[263:260] ^ 0);
  assign w91[13] = |(datain[259:256] ^ 5);
  assign w91[14] = |(datain[255:252] ^ 11);
  assign w91[15] = |(datain[251:248] ^ 9);
  assign w91[16] = |(datain[247:244] ^ 0);
  assign w91[17] = |(datain[243:240] ^ 0);
  assign w91[18] = |(datain[239:236] ^ 1);
  assign w91[19] = |(datain[235:232] ^ 2);
  assign w91[20] = |(datain[231:228] ^ 11);
  assign w91[21] = |(datain[227:224] ^ 10);
  assign w91[22] = |(datain[223:220] ^ 15);
  assign w91[23] = |(datain[219:216] ^ 1);
  assign w91[24] = |(datain[215:212] ^ 1);
  assign w91[25] = |(datain[211:208] ^ 2);
  assign w91[26] = |(datain[207:204] ^ 11);
  assign w91[27] = |(datain[203:200] ^ 4);
  assign w91[28] = |(datain[199:196] ^ 4);
  assign w91[29] = |(datain[195:192] ^ 0);
  assign w91[30] = |(datain[191:188] ^ 12);
  assign w91[31] = |(datain[187:184] ^ 13);
  assign w91[32] = |(datain[183:180] ^ 2);
  assign w91[33] = |(datain[179:176] ^ 1);
  assign w91[34] = |(datain[175:172] ^ 14);
  assign w91[35] = |(datain[171:168] ^ 8);
  assign w91[36] = |(datain[167:164] ^ 15);
  assign w91[37] = |(datain[163:160] ^ 7);
  assign w91[38] = |(datain[159:156] ^ 0);
  assign w91[39] = |(datain[155:152] ^ 4);
  assign w91[40] = |(datain[151:148] ^ 11);
  assign w91[41] = |(datain[147:144] ^ 4);
  assign w91[42] = |(datain[143:140] ^ 4);
  assign w91[43] = |(datain[139:136] ^ 0);
  assign w91[44] = |(datain[135:132] ^ 11);
  assign w91[45] = |(datain[131:128] ^ 9);
  assign w91[46] = |(datain[127:124] ^ 0);
  assign w91[47] = |(datain[123:120] ^ 3);
  assign w91[48] = |(datain[119:116] ^ 0);
  assign w91[49] = |(datain[115:112] ^ 0);
  assign w91[50] = |(datain[111:108] ^ 11);
  assign w91[51] = |(datain[107:104] ^ 10);
  assign w91[52] = |(datain[103:100] ^ 2);
  assign w91[53] = |(datain[99:96] ^ 9);
  assign w91[54] = |(datain[95:92] ^ 0);
  assign w91[55] = |(datain[91:88] ^ 11);
  assign w91[56] = |(datain[87:84] ^ 12);
  assign w91[57] = |(datain[83:80] ^ 13);
  assign w91[58] = |(datain[79:76] ^ 2);
  assign w91[59] = |(datain[75:72] ^ 1);
  assign w91[60] = |(datain[71:68] ^ 14);
  assign w91[61] = |(datain[67:64] ^ 9);
  assign w91[62] = |(datain[63:60] ^ 13);
  assign w91[63] = |(datain[59:56] ^ 7);
  assign w91[64] = |(datain[55:52] ^ 0);
  assign w91[65] = |(datain[51:48] ^ 0);
  assign w91[66] = |(datain[47:44] ^ 8);
  assign w91[67] = |(datain[43:40] ^ 0);
  assign w91[68] = |(datain[39:36] ^ 3);
  assign w91[69] = |(datain[35:32] ^ 14);
  assign w91[70] = |(datain[31:28] ^ 8);
  assign w91[71] = |(datain[27:24] ^ 2);
  assign w91[72] = |(datain[23:20] ^ 0);
  assign w91[73] = |(datain[19:16] ^ 11);
  assign comp[91] = ~(|w91);
  wire [76-1:0] w92;
  assign w92[0] = |(datain[311:308] ^ 11);
  assign w92[1] = |(datain[307:304] ^ 8);
  assign w92[2] = |(datain[303:300] ^ 0);
  assign w92[3] = |(datain[299:296] ^ 0);
  assign w92[4] = |(datain[295:292] ^ 4);
  assign w92[5] = |(datain[291:288] ^ 2);
  assign w92[6] = |(datain[287:284] ^ 3);
  assign w92[7] = |(datain[283:280] ^ 3);
  assign w92[8] = |(datain[279:276] ^ 12);
  assign w92[9] = |(datain[275:272] ^ 9);
  assign w92[10] = |(datain[271:268] ^ 3);
  assign w92[11] = |(datain[267:264] ^ 3);
  assign w92[12] = |(datain[263:260] ^ 13);
  assign w92[13] = |(datain[259:256] ^ 2);
  assign w92[14] = |(datain[255:252] ^ 12);
  assign w92[15] = |(datain[251:248] ^ 13);
  assign w92[16] = |(datain[247:244] ^ 0);
  assign w92[17] = |(datain[243:240] ^ 1);
  assign w92[18] = |(datain[239:236] ^ 11);
  assign w92[19] = |(datain[235:232] ^ 4);
  assign w92[20] = |(datain[231:228] ^ 4);
  assign w92[21] = |(datain[227:224] ^ 0);
  assign w92[22] = |(datain[223:220] ^ 11);
  assign w92[23] = |(datain[219:216] ^ 10);
  assign w92[24] = |(datain[215:212] ^ 14);
  assign w92[25] = |(datain[211:208] ^ 7);
  assign w92[26] = |(datain[207:204] ^ 0);
  assign w92[27] = |(datain[203:200] ^ 4);
  assign w92[28] = |(datain[199:196] ^ 11);
  assign w92[29] = |(datain[195:192] ^ 9);
  assign w92[30] = |(datain[191:188] ^ 0);
  assign w92[31] = |(datain[187:184] ^ 3);
  assign w92[32] = |(datain[183:180] ^ 0);
  assign w92[33] = |(datain[179:176] ^ 0);
  assign w92[34] = |(datain[175:172] ^ 12);
  assign w92[35] = |(datain[171:168] ^ 12);
  assign w92[36] = |(datain[167:164] ^ 5);
  assign w92[37] = |(datain[163:160] ^ 10);
  assign w92[38] = |(datain[159:156] ^ 5);
  assign w92[39] = |(datain[155:152] ^ 9);
  assign w92[40] = |(datain[151:148] ^ 11);
  assign w92[41] = |(datain[147:144] ^ 8);
  assign w92[42] = |(datain[143:140] ^ 0);
  assign w92[43] = |(datain[139:136] ^ 1);
  assign w92[44] = |(datain[135:132] ^ 5);
  assign w92[45] = |(datain[131:128] ^ 7);
  assign w92[46] = |(datain[127:124] ^ 12);
  assign w92[47] = |(datain[123:120] ^ 13);
  assign w92[48] = |(datain[119:116] ^ 0);
  assign w92[49] = |(datain[115:112] ^ 1);
  assign w92[50] = |(datain[111:108] ^ 11);
  assign w92[51] = |(datain[107:104] ^ 4);
  assign w92[52] = |(datain[103:100] ^ 3);
  assign w92[53] = |(datain[99:96] ^ 14);
  assign w92[54] = |(datain[95:92] ^ 12);
  assign w92[55] = |(datain[91:88] ^ 12);
  assign w92[56] = |(datain[87:84] ^ 11);
  assign w92[57] = |(datain[83:80] ^ 8);
  assign w92[58] = |(datain[79:76] ^ 0);
  assign w92[59] = |(datain[75:72] ^ 1);
  assign w92[60] = |(datain[71:68] ^ 4);
  assign w92[61] = |(datain[67:64] ^ 3);
  assign w92[62] = |(datain[63:60] ^ 5);
  assign w92[63] = |(datain[59:56] ^ 10);
  assign w92[64] = |(datain[55:52] ^ 1);
  assign w92[65] = |(datain[51:48] ^ 15);
  assign w92[66] = |(datain[47:44] ^ 5);
  assign w92[67] = |(datain[43:40] ^ 9);
  assign w92[68] = |(datain[39:36] ^ 12);
  assign w92[69] = |(datain[35:32] ^ 12);
  assign w92[70] = |(datain[31:28] ^ 14);
  assign w92[71] = |(datain[27:24] ^ 9);
  assign w92[72] = |(datain[23:20] ^ 13);
  assign w92[73] = |(datain[19:16] ^ 11);
  assign w92[74] = |(datain[15:12] ^ 15);
  assign w92[75] = |(datain[11:8] ^ 14);
  assign comp[92] = ~(|w92);
  wire [74-1:0] w93;
  assign w93[0] = |(datain[311:308] ^ 0);
  assign w93[1] = |(datain[307:304] ^ 8);
  assign w93[2] = |(datain[303:300] ^ 8);
  assign w93[3] = |(datain[299:296] ^ 1);
  assign w93[4] = |(datain[295:292] ^ 15);
  assign w93[5] = |(datain[291:288] ^ 11);
  assign w93[6] = |(datain[287:284] ^ 5);
  assign w93[7] = |(datain[283:280] ^ 3);
  assign w93[8] = |(datain[279:276] ^ 4);
  assign w93[9] = |(datain[275:272] ^ 2);
  assign w93[10] = |(datain[271:268] ^ 7);
  assign w93[11] = |(datain[267:264] ^ 5);
  assign w93[12] = |(datain[263:260] ^ 0);
  assign w93[13] = |(datain[259:256] ^ 2);
  assign w93[14] = |(datain[255:252] ^ 15);
  assign w93[15] = |(datain[251:248] ^ 9);
  assign w93[16] = |(datain[247:244] ^ 12);
  assign w93[17] = |(datain[243:240] ^ 3);
  assign w93[18] = |(datain[239:236] ^ 15);
  assign w93[19] = |(datain[235:232] ^ 8);
  assign w93[20] = |(datain[231:228] ^ 12);
  assign w93[21] = |(datain[227:224] ^ 3);
  assign w93[22] = |(datain[223:220] ^ 9);
  assign w93[23] = |(datain[219:216] ^ 12);
  assign w93[24] = |(datain[215:212] ^ 2);
  assign w93[25] = |(datain[211:208] ^ 14);
  assign w93[26] = |(datain[207:204] ^ 15);
  assign w93[27] = |(datain[203:200] ^ 15);
  assign w93[28] = |(datain[199:196] ^ 1);
  assign w93[29] = |(datain[195:192] ^ 14);
  assign w93[30] = |(datain[191:188] ^ 9);
  assign w93[31] = |(datain[187:184] ^ 0);
  assign w93[32] = |(datain[183:180] ^ 0);
  assign w93[33] = |(datain[179:176] ^ 6);
  assign w93[34] = |(datain[175:172] ^ 12);
  assign w93[35] = |(datain[171:168] ^ 3);
  assign w93[36] = |(datain[167:164] ^ 11);
  assign w93[37] = |(datain[163:160] ^ 0);
  assign w93[38] = |(datain[159:156] ^ 0);
  assign w93[39] = |(datain[155:152] ^ 3);
  assign w93[40] = |(datain[151:148] ^ 12);
  assign w93[41] = |(datain[147:144] ^ 15);
  assign w93[42] = |(datain[143:140] ^ 1);
  assign w93[43] = |(datain[139:136] ^ 14);
  assign w93[44] = |(datain[135:132] ^ 0);
  assign w93[45] = |(datain[131:128] ^ 6);
  assign w93[46] = |(datain[127:124] ^ 3);
  assign w93[47] = |(datain[123:120] ^ 3);
  assign w93[48] = |(datain[119:116] ^ 12);
  assign w93[49] = |(datain[115:112] ^ 0);
  assign w93[50] = |(datain[111:108] ^ 8);
  assign w93[51] = |(datain[107:104] ^ 14);
  assign w93[52] = |(datain[103:100] ^ 13);
  assign w93[53] = |(datain[99:96] ^ 8);
  assign w93[54] = |(datain[95:92] ^ 8);
  assign w93[55] = |(datain[91:88] ^ 12);
  assign w93[56] = |(datain[87:84] ^ 12);
  assign w93[57] = |(datain[83:80] ^ 8);
  assign w93[58] = |(datain[79:76] ^ 8);
  assign w93[59] = |(datain[75:72] ^ 14);
  assign w93[60] = |(datain[71:68] ^ 12);
  assign w93[61] = |(datain[67:64] ^ 0);
  assign w93[62] = |(datain[63:60] ^ 11);
  assign w93[63] = |(datain[59:56] ^ 14);
  assign w93[64] = |(datain[55:52] ^ 9);
  assign w93[65] = |(datain[51:48] ^ 0);
  assign w93[66] = |(datain[47:44] ^ 0);
  assign w93[67] = |(datain[43:40] ^ 0);
  assign w93[68] = |(datain[39:36] ^ 11);
  assign w93[69] = |(datain[35:32] ^ 15);
  assign w93[70] = |(datain[31:28] ^ 15);
  assign w93[71] = |(datain[27:24] ^ 11);
  assign w93[72] = |(datain[23:20] ^ 0);
  assign w93[73] = |(datain[19:16] ^ 5);
  assign comp[93] = ~(|w93);
  wire [76-1:0] w94;
  assign w94[0] = |(datain[311:308] ^ 2);
  assign w94[1] = |(datain[307:304] ^ 13);
  assign w94[2] = |(datain[303:300] ^ 0);
  assign w94[3] = |(datain[299:296] ^ 3);
  assign w94[4] = |(datain[295:292] ^ 0);
  assign w94[5] = |(datain[291:288] ^ 0);
  assign w94[6] = |(datain[287:284] ^ 8);
  assign w94[7] = |(datain[283:280] ^ 9);
  assign w94[8] = |(datain[279:276] ^ 8);
  assign w94[9] = |(datain[275:272] ^ 6);
  assign w94[10] = |(datain[271:268] ^ 11);
  assign w94[11] = |(datain[267:264] ^ 9);
  assign w94[12] = |(datain[263:260] ^ 0);
  assign w94[13] = |(datain[259:256] ^ 0);
  assign w94[14] = |(datain[255:252] ^ 11);
  assign w94[15] = |(datain[251:248] ^ 4);
  assign w94[16] = |(datain[247:244] ^ 4);
  assign w94[17] = |(datain[243:240] ^ 0);
  assign w94[18] = |(datain[239:236] ^ 11);
  assign w94[19] = |(datain[235:232] ^ 9);
  assign w94[20] = |(datain[231:228] ^ 11);
  assign w94[21] = |(datain[227:224] ^ 6);
  assign w94[22] = |(datain[223:220] ^ 0);
  assign w94[23] = |(datain[219:216] ^ 0);
  assign w94[24] = |(datain[215:212] ^ 8);
  assign w94[25] = |(datain[211:208] ^ 13);
  assign w94[26] = |(datain[207:204] ^ 9);
  assign w94[27] = |(datain[203:200] ^ 6);
  assign w94[28] = |(datain[199:196] ^ 0);
  assign w94[29] = |(datain[195:192] ^ 3);
  assign w94[30] = |(datain[191:188] ^ 0);
  assign w94[31] = |(datain[187:184] ^ 0);
  assign w94[32] = |(datain[183:180] ^ 12);
  assign w94[33] = |(datain[179:176] ^ 13);
  assign w94[34] = |(datain[175:172] ^ 2);
  assign w94[35] = |(datain[171:168] ^ 1);
  assign w94[36] = |(datain[167:164] ^ 11);
  assign w94[37] = |(datain[163:160] ^ 0);
  assign w94[38] = |(datain[159:156] ^ 0);
  assign w94[39] = |(datain[155:152] ^ 0);
  assign w94[40] = |(datain[151:148] ^ 14);
  assign w94[41] = |(datain[147:144] ^ 8);
  assign w94[42] = |(datain[143:140] ^ 1);
  assign w94[43] = |(datain[139:136] ^ 11);
  assign w94[44] = |(datain[135:132] ^ 0);
  assign w94[45] = |(datain[131:128] ^ 0);
  assign w94[46] = |(datain[127:124] ^ 11);
  assign w94[47] = |(datain[123:120] ^ 4);
  assign w94[48] = |(datain[119:116] ^ 4);
  assign w94[49] = |(datain[115:112] ^ 0);
  assign w94[50] = |(datain[111:108] ^ 11);
  assign w94[51] = |(datain[107:104] ^ 9);
  assign w94[52] = |(datain[103:100] ^ 0);
  assign w94[53] = |(datain[99:96] ^ 3);
  assign w94[54] = |(datain[95:92] ^ 0);
  assign w94[55] = |(datain[91:88] ^ 0);
  assign w94[56] = |(datain[87:84] ^ 8);
  assign w94[57] = |(datain[83:80] ^ 13);
  assign w94[58] = |(datain[79:76] ^ 9);
  assign w94[59] = |(datain[75:72] ^ 6);
  assign w94[60] = |(datain[71:68] ^ 11);
  assign w94[61] = |(datain[67:64] ^ 8);
  assign w94[62] = |(datain[63:60] ^ 0);
  assign w94[63] = |(datain[59:56] ^ 0);
  assign w94[64] = |(datain[55:52] ^ 12);
  assign w94[65] = |(datain[51:48] ^ 13);
  assign w94[66] = |(datain[47:44] ^ 2);
  assign w94[67] = |(datain[43:40] ^ 1);
  assign w94[68] = |(datain[39:36] ^ 5);
  assign w94[69] = |(datain[35:32] ^ 10);
  assign w94[70] = |(datain[31:28] ^ 5);
  assign w94[71] = |(datain[27:24] ^ 9);
  assign w94[72] = |(datain[23:20] ^ 8);
  assign w94[73] = |(datain[19:16] ^ 3);
  assign w94[74] = |(datain[15:12] ^ 12);
  assign w94[75] = |(datain[11:8] ^ 9);
  assign comp[94] = ~(|w94);
  wire [76-1:0] w95;
  assign w95[0] = |(datain[311:308] ^ 2);
  assign w95[1] = |(datain[307:304] ^ 13);
  assign w95[2] = |(datain[303:300] ^ 0);
  assign w95[3] = |(datain[299:296] ^ 3);
  assign w95[4] = |(datain[295:292] ^ 0);
  assign w95[5] = |(datain[291:288] ^ 0);
  assign w95[6] = |(datain[287:284] ^ 8);
  assign w95[7] = |(datain[283:280] ^ 9);
  assign w95[8] = |(datain[279:276] ^ 8);
  assign w95[9] = |(datain[275:272] ^ 6);
  assign w95[10] = |(datain[271:268] ^ 11);
  assign w95[11] = |(datain[267:264] ^ 11);
  assign w95[12] = |(datain[263:260] ^ 0);
  assign w95[13] = |(datain[259:256] ^ 0);
  assign w95[14] = |(datain[255:252] ^ 11);
  assign w95[15] = |(datain[251:248] ^ 4);
  assign w95[16] = |(datain[247:244] ^ 4);
  assign w95[17] = |(datain[243:240] ^ 0);
  assign w95[18] = |(datain[239:236] ^ 11);
  assign w95[19] = |(datain[235:232] ^ 9);
  assign w95[20] = |(datain[231:228] ^ 11);
  assign w95[21] = |(datain[227:224] ^ 8);
  assign w95[22] = |(datain[223:220] ^ 0);
  assign w95[23] = |(datain[219:216] ^ 0);
  assign w95[24] = |(datain[215:212] ^ 8);
  assign w95[25] = |(datain[211:208] ^ 13);
  assign w95[26] = |(datain[207:204] ^ 9);
  assign w95[27] = |(datain[203:200] ^ 6);
  assign w95[28] = |(datain[199:196] ^ 0);
  assign w95[29] = |(datain[195:192] ^ 3);
  assign w95[30] = |(datain[191:188] ^ 0);
  assign w95[31] = |(datain[187:184] ^ 0);
  assign w95[32] = |(datain[183:180] ^ 12);
  assign w95[33] = |(datain[179:176] ^ 13);
  assign w95[34] = |(datain[175:172] ^ 2);
  assign w95[35] = |(datain[171:168] ^ 1);
  assign w95[36] = |(datain[167:164] ^ 11);
  assign w95[37] = |(datain[163:160] ^ 0);
  assign w95[38] = |(datain[159:156] ^ 0);
  assign w95[39] = |(datain[155:152] ^ 0);
  assign w95[40] = |(datain[151:148] ^ 14);
  assign w95[41] = |(datain[147:144] ^ 8);
  assign w95[42] = |(datain[143:140] ^ 1);
  assign w95[43] = |(datain[139:136] ^ 11);
  assign w95[44] = |(datain[135:132] ^ 0);
  assign w95[45] = |(datain[131:128] ^ 0);
  assign w95[46] = |(datain[127:124] ^ 11);
  assign w95[47] = |(datain[123:120] ^ 4);
  assign w95[48] = |(datain[119:116] ^ 4);
  assign w95[49] = |(datain[115:112] ^ 0);
  assign w95[50] = |(datain[111:108] ^ 11);
  assign w95[51] = |(datain[107:104] ^ 9);
  assign w95[52] = |(datain[103:100] ^ 0);
  assign w95[53] = |(datain[99:96] ^ 3);
  assign w95[54] = |(datain[95:92] ^ 0);
  assign w95[55] = |(datain[91:88] ^ 0);
  assign w95[56] = |(datain[87:84] ^ 8);
  assign w95[57] = |(datain[83:80] ^ 13);
  assign w95[58] = |(datain[79:76] ^ 9);
  assign w95[59] = |(datain[75:72] ^ 6);
  assign w95[60] = |(datain[71:68] ^ 11);
  assign w95[61] = |(datain[67:64] ^ 10);
  assign w95[62] = |(datain[63:60] ^ 0);
  assign w95[63] = |(datain[59:56] ^ 0);
  assign w95[64] = |(datain[55:52] ^ 12);
  assign w95[65] = |(datain[51:48] ^ 13);
  assign w95[66] = |(datain[47:44] ^ 2);
  assign w95[67] = |(datain[43:40] ^ 1);
  assign w95[68] = |(datain[39:36] ^ 5);
  assign w95[69] = |(datain[35:32] ^ 10);
  assign w95[70] = |(datain[31:28] ^ 5);
  assign w95[71] = |(datain[27:24] ^ 9);
  assign w95[72] = |(datain[23:20] ^ 8);
  assign w95[73] = |(datain[19:16] ^ 3);
  assign w95[74] = |(datain[15:12] ^ 12);
  assign w95[75] = |(datain[11:8] ^ 9);
  assign comp[95] = ~(|w95);
  wire [76-1:0] w96;
  assign w96[0] = |(datain[311:308] ^ 12);
  assign w96[1] = |(datain[307:304] ^ 13);
  assign w96[2] = |(datain[303:300] ^ 2);
  assign w96[3] = |(datain[299:296] ^ 1);
  assign w96[4] = |(datain[295:292] ^ 11);
  assign w96[5] = |(datain[291:288] ^ 0);
  assign w96[6] = |(datain[287:284] ^ 0);
  assign w96[7] = |(datain[283:280] ^ 0);
  assign w96[8] = |(datain[279:276] ^ 14);
  assign w96[9] = |(datain[275:272] ^ 8);
  assign w96[10] = |(datain[271:268] ^ 1);
  assign w96[11] = |(datain[267:264] ^ 11);
  assign w96[12] = |(datain[263:260] ^ 0);
  assign w96[13] = |(datain[259:256] ^ 0);
  assign w96[14] = |(datain[255:252] ^ 11);
  assign w96[15] = |(datain[251:248] ^ 4);
  assign w96[16] = |(datain[247:244] ^ 4);
  assign w96[17] = |(datain[243:240] ^ 0);
  assign w96[18] = |(datain[239:236] ^ 11);
  assign w96[19] = |(datain[235:232] ^ 9);
  assign w96[20] = |(datain[231:228] ^ 0);
  assign w96[21] = |(datain[227:224] ^ 3);
  assign w96[22] = |(datain[223:220] ^ 0);
  assign w96[23] = |(datain[219:216] ^ 0);
  assign w96[24] = |(datain[215:212] ^ 8);
  assign w96[25] = |(datain[211:208] ^ 13);
  assign w96[26] = |(datain[207:204] ^ 9);
  assign w96[27] = |(datain[203:200] ^ 6);
  assign w96[28] = |(datain[199:196] ^ 11);
  assign w96[29] = |(datain[195:192] ^ 10);
  assign w96[30] = |(datain[191:188] ^ 0);
  assign w96[31] = |(datain[187:184] ^ 0);
  assign w96[32] = |(datain[183:180] ^ 12);
  assign w96[33] = |(datain[179:176] ^ 13);
  assign w96[34] = |(datain[175:172] ^ 2);
  assign w96[35] = |(datain[171:168] ^ 1);
  assign w96[36] = |(datain[167:164] ^ 5);
  assign w96[37] = |(datain[163:160] ^ 10);
  assign w96[38] = |(datain[159:156] ^ 5);
  assign w96[39] = |(datain[155:152] ^ 9);
  assign w96[40] = |(datain[151:148] ^ 8);
  assign w96[41] = |(datain[147:144] ^ 3);
  assign w96[42] = |(datain[143:140] ^ 12);
  assign w96[43] = |(datain[139:136] ^ 9);
  assign w96[44] = |(datain[135:132] ^ 1);
  assign w96[45] = |(datain[131:128] ^ 15);
  assign w96[46] = |(datain[127:124] ^ 11);
  assign w96[47] = |(datain[123:120] ^ 8);
  assign w96[48] = |(datain[119:116] ^ 0);
  assign w96[49] = |(datain[115:112] ^ 1);
  assign w96[50] = |(datain[111:108] ^ 5);
  assign w96[51] = |(datain[107:104] ^ 7);
  assign w96[52] = |(datain[103:100] ^ 12);
  assign w96[53] = |(datain[99:96] ^ 13);
  assign w96[54] = |(datain[95:92] ^ 2);
  assign w96[55] = |(datain[91:88] ^ 1);
  assign w96[56] = |(datain[87:84] ^ 11);
  assign w96[57] = |(datain[83:80] ^ 4);
  assign w96[58] = |(datain[79:76] ^ 3);
  assign w96[59] = |(datain[75:72] ^ 14);
  assign w96[60] = |(datain[71:68] ^ 12);
  assign w96[61] = |(datain[67:64] ^ 13);
  assign w96[62] = |(datain[63:60] ^ 2);
  assign w96[63] = |(datain[59:56] ^ 1);
  assign w96[64] = |(datain[55:52] ^ 14);
  assign w96[65] = |(datain[51:48] ^ 11);
  assign w96[66] = |(datain[47:44] ^ 8);
  assign w96[67] = |(datain[43:40] ^ 11);
  assign w96[68] = |(datain[39:36] ^ 3);
  assign w96[69] = |(datain[35:32] ^ 3);
  assign w96[70] = |(datain[31:28] ^ 12);
  assign w96[71] = |(datain[27:24] ^ 9);
  assign w96[72] = |(datain[23:20] ^ 3);
  assign w96[73] = |(datain[19:16] ^ 3);
  assign w96[74] = |(datain[15:12] ^ 13);
  assign w96[75] = |(datain[11:8] ^ 2);
  assign comp[96] = ~(|w96);
  wire [74-1:0] w97;
  assign w97[0] = |(datain[311:308] ^ 2);
  assign w97[1] = |(datain[307:304] ^ 1);
  assign w97[2] = |(datain[303:300] ^ 11);
  assign w97[3] = |(datain[299:296] ^ 0);
  assign w97[4] = |(datain[295:292] ^ 0);
  assign w97[5] = |(datain[291:288] ^ 0);
  assign w97[6] = |(datain[287:284] ^ 14);
  assign w97[7] = |(datain[283:280] ^ 8);
  assign w97[8] = |(datain[279:276] ^ 1);
  assign w97[9] = |(datain[275:272] ^ 12);
  assign w97[10] = |(datain[271:268] ^ 0);
  assign w97[11] = |(datain[267:264] ^ 0);
  assign w97[12] = |(datain[263:260] ^ 11);
  assign w97[13] = |(datain[259:256] ^ 4);
  assign w97[14] = |(datain[255:252] ^ 4);
  assign w97[15] = |(datain[251:248] ^ 0);
  assign w97[16] = |(datain[247:244] ^ 11);
  assign w97[17] = |(datain[243:240] ^ 9);
  assign w97[18] = |(datain[239:236] ^ 0);
  assign w97[19] = |(datain[235:232] ^ 3);
  assign w97[20] = |(datain[231:228] ^ 0);
  assign w97[21] = |(datain[227:224] ^ 0);
  assign w97[22] = |(datain[223:220] ^ 8);
  assign w97[23] = |(datain[219:216] ^ 13);
  assign w97[24] = |(datain[215:212] ^ 9);
  assign w97[25] = |(datain[211:208] ^ 6);
  assign w97[26] = |(datain[207:204] ^ 12);
  assign w97[27] = |(datain[203:200] ^ 15);
  assign w97[28] = |(datain[199:196] ^ 0);
  assign w97[29] = |(datain[195:192] ^ 0);
  assign w97[30] = |(datain[191:188] ^ 12);
  assign w97[31] = |(datain[187:184] ^ 13);
  assign w97[32] = |(datain[183:180] ^ 2);
  assign w97[33] = |(datain[179:176] ^ 1);
  assign w97[34] = |(datain[175:172] ^ 5);
  assign w97[35] = |(datain[171:168] ^ 10);
  assign w97[36] = |(datain[167:164] ^ 5);
  assign w97[37] = |(datain[163:160] ^ 9);
  assign w97[38] = |(datain[159:156] ^ 8);
  assign w97[39] = |(datain[155:152] ^ 3);
  assign w97[40] = |(datain[151:148] ^ 12);
  assign w97[41] = |(datain[147:144] ^ 9);
  assign w97[42] = |(datain[143:140] ^ 1);
  assign w97[43] = |(datain[139:136] ^ 15);
  assign w97[44] = |(datain[135:132] ^ 11);
  assign w97[45] = |(datain[131:128] ^ 8);
  assign w97[46] = |(datain[127:124] ^ 0);
  assign w97[47] = |(datain[123:120] ^ 1);
  assign w97[48] = |(datain[119:116] ^ 5);
  assign w97[49] = |(datain[115:112] ^ 7);
  assign w97[50] = |(datain[111:108] ^ 12);
  assign w97[51] = |(datain[107:104] ^ 13);
  assign w97[52] = |(datain[103:100] ^ 2);
  assign w97[53] = |(datain[99:96] ^ 1);
  assign w97[54] = |(datain[95:92] ^ 11);
  assign w97[55] = |(datain[91:88] ^ 4);
  assign w97[56] = |(datain[87:84] ^ 3);
  assign w97[57] = |(datain[83:80] ^ 14);
  assign w97[58] = |(datain[79:76] ^ 12);
  assign w97[59] = |(datain[75:72] ^ 13);
  assign w97[60] = |(datain[71:68] ^ 2);
  assign w97[61] = |(datain[67:64] ^ 1);
  assign w97[62] = |(datain[63:60] ^ 14);
  assign w97[63] = |(datain[59:56] ^ 9);
  assign w97[64] = |(datain[55:52] ^ 7);
  assign w97[65] = |(datain[51:48] ^ 6);
  assign w97[66] = |(datain[47:44] ^ 15);
  assign w97[67] = |(datain[43:40] ^ 15);
  assign w97[68] = |(datain[39:36] ^ 3);
  assign w97[69] = |(datain[35:32] ^ 3);
  assign w97[70] = |(datain[31:28] ^ 12);
  assign w97[71] = |(datain[27:24] ^ 9);
  assign w97[72] = |(datain[23:20] ^ 3);
  assign w97[73] = |(datain[19:16] ^ 3);
  assign comp[97] = ~(|w97);
  wire [76-1:0] w98;
  assign w98[0] = |(datain[311:308] ^ 0);
  assign w98[1] = |(datain[307:304] ^ 2);
  assign w98[2] = |(datain[303:300] ^ 3);
  assign w98[3] = |(datain[299:296] ^ 13);
  assign w98[4] = |(datain[295:292] ^ 11);
  assign w98[5] = |(datain[291:288] ^ 10);
  assign w98[6] = |(datain[287:284] ^ 9);
  assign w98[7] = |(datain[283:280] ^ 14);
  assign w98[8] = |(datain[279:276] ^ 0);
  assign w98[9] = |(datain[275:272] ^ 0);
  assign w98[10] = |(datain[271:268] ^ 12);
  assign w98[11] = |(datain[267:264] ^ 13);
  assign w98[12] = |(datain[263:260] ^ 2);
  assign w98[13] = |(datain[259:256] ^ 1);
  assign w98[14] = |(datain[255:252] ^ 9);
  assign w98[15] = |(datain[251:248] ^ 3);
  assign w98[16] = |(datain[247:244] ^ 11);
  assign w98[17] = |(datain[243:240] ^ 4);
  assign w98[18] = |(datain[239:236] ^ 4);
  assign w98[19] = |(datain[235:232] ^ 0);
  assign w98[20] = |(datain[231:228] ^ 11);
  assign w98[21] = |(datain[227:224] ^ 9);
  assign w98[22] = |(datain[223:220] ^ 11);
  assign w98[23] = |(datain[219:216] ^ 4);
  assign w98[24] = |(datain[215:212] ^ 0);
  assign w98[25] = |(datain[211:208] ^ 0);
  assign w98[26] = |(datain[207:204] ^ 11);
  assign w98[27] = |(datain[203:200] ^ 10);
  assign w98[28] = |(datain[199:196] ^ 0);
  assign w98[29] = |(datain[195:192] ^ 0);
  assign w98[30] = |(datain[191:188] ^ 0);
  assign w98[31] = |(datain[187:184] ^ 1);
  assign w98[32] = |(datain[183:180] ^ 12);
  assign w98[33] = |(datain[179:176] ^ 13);
  assign w98[34] = |(datain[175:172] ^ 2);
  assign w98[35] = |(datain[171:168] ^ 1);
  assign w98[36] = |(datain[167:164] ^ 11);
  assign w98[37] = |(datain[163:160] ^ 4);
  assign w98[38] = |(datain[159:156] ^ 3);
  assign w98[39] = |(datain[155:152] ^ 14);
  assign w98[40] = |(datain[151:148] ^ 12);
  assign w98[41] = |(datain[147:144] ^ 13);
  assign w98[42] = |(datain[143:140] ^ 2);
  assign w98[43] = |(datain[139:136] ^ 1);
  assign w98[44] = |(datain[135:132] ^ 11);
  assign w98[45] = |(datain[131:128] ^ 4);
  assign w98[46] = |(datain[127:124] ^ 4);
  assign w98[47] = |(datain[123:120] ^ 15);
  assign w98[48] = |(datain[119:116] ^ 14);
  assign w98[49] = |(datain[115:112] ^ 11);
  assign w98[50] = |(datain[111:108] ^ 13);
  assign w98[51] = |(datain[107:104] ^ 12);
  assign w98[52] = |(datain[103:100] ^ 11);
  assign w98[53] = |(datain[99:96] ^ 4);
  assign w98[54] = |(datain[95:92] ^ 0);
  assign w98[55] = |(datain[91:88] ^ 9);
  assign w98[56] = |(datain[87:84] ^ 11);
  assign w98[57] = |(datain[83:80] ^ 10);
  assign w98[58] = |(datain[79:76] ^ 3);
  assign w98[59] = |(datain[75:72] ^ 5);
  assign w98[60] = |(datain[71:68] ^ 0);
  assign w98[61] = |(datain[67:64] ^ 1);
  assign w98[62] = |(datain[63:60] ^ 12);
  assign w98[63] = |(datain[59:56] ^ 13);
  assign w98[64] = |(datain[55:52] ^ 2);
  assign w98[65] = |(datain[51:48] ^ 1);
  assign w98[66] = |(datain[47:44] ^ 12);
  assign w98[67] = |(datain[43:40] ^ 13);
  assign w98[68] = |(datain[39:36] ^ 2);
  assign w98[69] = |(datain[35:32] ^ 0);
  assign w98[70] = |(datain[31:28] ^ 2);
  assign w98[71] = |(datain[27:24] ^ 10);
  assign w98[72] = |(datain[23:20] ^ 2);
  assign w98[73] = |(datain[19:16] ^ 14);
  assign w98[74] = |(datain[15:12] ^ 6);
  assign w98[75] = |(datain[11:8] ^ 3);
  assign comp[98] = ~(|w98);
  wire [76-1:0] w99;
  assign w99[0] = |(datain[311:308] ^ 4);
  assign w99[1] = |(datain[307:304] ^ 2);
  assign w99[2] = |(datain[303:300] ^ 3);
  assign w99[3] = |(datain[299:296] ^ 3);
  assign w99[4] = |(datain[295:292] ^ 12);
  assign w99[5] = |(datain[291:288] ^ 9);
  assign w99[6] = |(datain[287:284] ^ 3);
  assign w99[7] = |(datain[283:280] ^ 3);
  assign w99[8] = |(datain[279:276] ^ 13);
  assign w99[9] = |(datain[275:272] ^ 2);
  assign w99[10] = |(datain[271:268] ^ 12);
  assign w99[11] = |(datain[267:264] ^ 13);
  assign w99[12] = |(datain[263:260] ^ 2);
  assign w99[13] = |(datain[259:256] ^ 1);
  assign w99[14] = |(datain[255:252] ^ 11);
  assign w99[15] = |(datain[251:248] ^ 4);
  assign w99[16] = |(datain[247:244] ^ 4);
  assign w99[17] = |(datain[243:240] ^ 0);
  assign w99[18] = |(datain[239:236] ^ 8);
  assign w99[19] = |(datain[235:232] ^ 13);
  assign w99[20] = |(datain[231:228] ^ 9);
  assign w99[21] = |(datain[227:224] ^ 6);
  assign w99[22] = |(datain[223:220] ^ 12);
  assign w99[23] = |(datain[219:216] ^ 15);
  assign w99[24] = |(datain[215:212] ^ 0);
  assign w99[25] = |(datain[211:208] ^ 2);
  assign w99[26] = |(datain[207:204] ^ 11);
  assign w99[27] = |(datain[203:200] ^ 9);
  assign w99[28] = |(datain[199:196] ^ 1);
  assign w99[29] = |(datain[195:192] ^ 10);
  assign w99[30] = |(datain[191:188] ^ 0);
  assign w99[31] = |(datain[187:184] ^ 0);
  assign w99[32] = |(datain[183:180] ^ 12);
  assign w99[33] = |(datain[179:176] ^ 13);
  assign w99[34] = |(datain[175:172] ^ 2);
  assign w99[35] = |(datain[171:168] ^ 1);
  assign w99[36] = |(datain[167:164] ^ 11);
  assign w99[37] = |(datain[163:160] ^ 4);
  assign w99[38] = |(datain[159:156] ^ 3);
  assign w99[39] = |(datain[155:152] ^ 14);
  assign w99[40] = |(datain[151:148] ^ 12);
  assign w99[41] = |(datain[147:144] ^ 13);
  assign w99[42] = |(datain[143:140] ^ 2);
  assign w99[43] = |(datain[139:136] ^ 1);
  assign w99[44] = |(datain[135:132] ^ 12);
  assign w99[45] = |(datain[131:128] ^ 3);
  assign w99[46] = |(datain[127:124] ^ 11);
  assign w99[47] = |(datain[123:120] ^ 0);
  assign w99[48] = |(datain[119:116] ^ 0);
  assign w99[49] = |(datain[115:112] ^ 3);
  assign w99[50] = |(datain[111:108] ^ 12);
  assign w99[51] = |(datain[107:104] ^ 15);
  assign w99[52] = |(datain[103:100] ^ 11);
  assign w99[53] = |(datain[99:96] ^ 8);
  assign w99[54] = |(datain[95:92] ^ 2);
  assign w99[55] = |(datain[91:88] ^ 4);
  assign w99[56] = |(datain[87:84] ^ 3);
  assign w99[57] = |(datain[83:80] ^ 5);
  assign w99[58] = |(datain[79:76] ^ 12);
  assign w99[59] = |(datain[75:72] ^ 13);
  assign w99[60] = |(datain[71:68] ^ 2);
  assign w99[61] = |(datain[67:64] ^ 1);
  assign w99[62] = |(datain[63:60] ^ 5);
  assign w99[63] = |(datain[59:56] ^ 3);
  assign w99[64] = |(datain[55:52] ^ 0);
  assign w99[65] = |(datain[51:48] ^ 6);
  assign w99[66] = |(datain[47:44] ^ 11);
  assign w99[67] = |(datain[43:40] ^ 4);
  assign w99[68] = |(datain[39:36] ^ 2);
  assign w99[69] = |(datain[35:32] ^ 5);
  assign w99[70] = |(datain[31:28] ^ 8);
  assign w99[71] = |(datain[27:24] ^ 13);
  assign w99[72] = |(datain[23:20] ^ 9);
  assign w99[73] = |(datain[19:16] ^ 6);
  assign w99[74] = |(datain[15:12] ^ 15);
  assign w99[75] = |(datain[11:8] ^ 0);
  assign comp[99] = ~(|w99);
  wire [76-1:0] w100;
  assign w100[0] = |(datain[311:308] ^ 0);
  assign w100[1] = |(datain[307:304] ^ 1);
  assign w100[2] = |(datain[303:300] ^ 8);
  assign w100[3] = |(datain[299:296] ^ 11);
  assign w100[4] = |(datain[295:292] ^ 1);
  assign w100[5] = |(datain[291:288] ^ 14);
  assign w100[6] = |(datain[287:284] ^ 10);
  assign w100[7] = |(datain[283:280] ^ 11);
  assign w100[8] = |(datain[279:276] ^ 0);
  assign w100[9] = |(datain[275:272] ^ 6);
  assign w100[10] = |(datain[271:268] ^ 14);
  assign w100[11] = |(datain[267:264] ^ 8);
  assign w100[12] = |(datain[263:260] ^ 1);
  assign w100[13] = |(datain[259:256] ^ 8);
  assign w100[14] = |(datain[255:252] ^ 0);
  assign w100[15] = |(datain[251:248] ^ 1);
  assign w100[16] = |(datain[247:244] ^ 11);
  assign w100[17] = |(datain[243:240] ^ 4);
  assign w100[18] = |(datain[239:236] ^ 4);
  assign w100[19] = |(datain[235:232] ^ 0);
  assign w100[20] = |(datain[231:228] ^ 11);
  assign w100[21] = |(datain[227:224] ^ 9);
  assign w100[22] = |(datain[223:220] ^ 10);
  assign w100[23] = |(datain[219:216] ^ 9);
  assign w100[24] = |(datain[215:212] ^ 0);
  assign w100[25] = |(datain[211:208] ^ 6);
  assign w100[26] = |(datain[207:204] ^ 11);
  assign w100[27] = |(datain[203:200] ^ 10);
  assign w100[28] = |(datain[199:196] ^ 11);
  assign w100[29] = |(datain[195:192] ^ 6);
  assign w100[30] = |(datain[191:188] ^ 0);
  assign w100[31] = |(datain[187:184] ^ 6);
  assign w100[32] = |(datain[183:180] ^ 12);
  assign w100[33] = |(datain[179:176] ^ 13);
  assign w100[34] = |(datain[175:172] ^ 2);
  assign w100[35] = |(datain[171:168] ^ 1);
  assign w100[36] = |(datain[167:164] ^ 2);
  assign w100[37] = |(datain[163:160] ^ 6);
  assign w100[38] = |(datain[159:156] ^ 12);
  assign w100[39] = |(datain[155:152] ^ 7);
  assign w100[40] = |(datain[151:148] ^ 4);
  assign w100[41] = |(datain[147:144] ^ 5);
  assign w100[42] = |(datain[143:140] ^ 1);
  assign w100[43] = |(datain[139:136] ^ 5);
  assign w100[44] = |(datain[135:132] ^ 0);
  assign w100[45] = |(datain[131:128] ^ 0);
  assign w100[46] = |(datain[127:124] ^ 0);
  assign w100[47] = |(datain[123:120] ^ 0);
  assign w100[48] = |(datain[119:116] ^ 2);
  assign w100[49] = |(datain[115:112] ^ 6);
  assign w100[50] = |(datain[111:108] ^ 12);
  assign w100[51] = |(datain[107:104] ^ 7);
  assign w100[52] = |(datain[103:100] ^ 4);
  assign w100[53] = |(datain[99:96] ^ 5);
  assign w100[54] = |(datain[95:92] ^ 1);
  assign w100[55] = |(datain[91:88] ^ 7);
  assign w100[56] = |(datain[87:84] ^ 0);
  assign w100[57] = |(datain[83:80] ^ 0);
  assign w100[58] = |(datain[79:76] ^ 0);
  assign w100[59] = |(datain[75:72] ^ 0);
  assign w100[60] = |(datain[71:68] ^ 11);
  assign w100[61] = |(datain[67:64] ^ 4);
  assign w100[62] = |(datain[63:60] ^ 4);
  assign w100[63] = |(datain[59:56] ^ 0);
  assign w100[64] = |(datain[55:52] ^ 11);
  assign w100[65] = |(datain[51:48] ^ 9);
  assign w100[66] = |(datain[47:44] ^ 0);
  assign w100[67] = |(datain[43:40] ^ 3);
  assign w100[68] = |(datain[39:36] ^ 0);
  assign w100[69] = |(datain[35:32] ^ 0);
  assign w100[70] = |(datain[31:28] ^ 11);
  assign w100[71] = |(datain[27:24] ^ 10);
  assign w100[72] = |(datain[23:20] ^ 7);
  assign w100[73] = |(datain[19:16] ^ 10);
  assign w100[74] = |(datain[15:12] ^ 0);
  assign w100[75] = |(datain[11:8] ^ 6);
  assign comp[100] = ~(|w100);
  wire [74-1:0] w101;
  assign w101[0] = |(datain[311:308] ^ 0);
  assign w101[1] = |(datain[307:304] ^ 2);
  assign w101[2] = |(datain[303:300] ^ 11);
  assign w101[3] = |(datain[299:296] ^ 10);
  assign w101[4] = |(datain[295:292] ^ 0);
  assign w101[5] = |(datain[291:288] ^ 3);
  assign w101[6] = |(datain[287:284] ^ 0);
  assign w101[7] = |(datain[283:280] ^ 1);
  assign w101[8] = |(datain[279:276] ^ 0);
  assign w101[9] = |(datain[275:272] ^ 3);
  assign w101[10] = |(datain[271:268] ^ 1);
  assign w101[11] = |(datain[267:264] ^ 6);
  assign w101[12] = |(datain[263:260] ^ 0);
  assign w101[13] = |(datain[259:256] ^ 6);
  assign w101[14] = |(datain[255:252] ^ 0);
  assign w101[15] = |(datain[251:248] ^ 1);
  assign w101[16] = |(datain[247:244] ^ 8);
  assign w101[17] = |(datain[243:240] ^ 3);
  assign w101[18] = |(datain[239:236] ^ 14);
  assign w101[19] = |(datain[235:232] ^ 10);
  assign w101[20] = |(datain[231:228] ^ 0);
  assign w101[21] = |(datain[227:224] ^ 3);
  assign w101[22] = |(datain[223:220] ^ 2);
  assign w101[23] = |(datain[219:216] ^ 11);
  assign w101[24] = |(datain[215:212] ^ 12);
  assign w101[25] = |(datain[211:208] ^ 10);
  assign w101[26] = |(datain[207:204] ^ 11);
  assign w101[27] = |(datain[203:200] ^ 4);
  assign w101[28] = |(datain[199:196] ^ 4);
  assign w101[29] = |(datain[195:192] ^ 0);
  assign w101[30] = |(datain[191:188] ^ 12);
  assign w101[31] = |(datain[187:184] ^ 13);
  assign w101[32] = |(datain[183:180] ^ 2);
  assign w101[33] = |(datain[179:176] ^ 1);
  assign w101[34] = |(datain[175:172] ^ 7);
  assign w101[35] = |(datain[171:168] ^ 2);
  assign w101[36] = |(datain[167:164] ^ 1);
  assign w101[37] = |(datain[163:160] ^ 4);
  assign w101[38] = |(datain[159:156] ^ 9);
  assign w101[39] = |(datain[155:152] ^ 0);
  assign w101[40] = |(datain[151:148] ^ 9);
  assign w101[41] = |(datain[147:144] ^ 0);
  assign w101[42] = |(datain[143:140] ^ 9);
  assign w101[43] = |(datain[139:136] ^ 0);
  assign w101[44] = |(datain[135:132] ^ 11);
  assign w101[45] = |(datain[131:128] ^ 8);
  assign w101[46] = |(datain[127:124] ^ 0);
  assign w101[47] = |(datain[123:120] ^ 0);
  assign w101[48] = |(datain[119:116] ^ 5);
  assign w101[49] = |(datain[115:112] ^ 7);
  assign w101[50] = |(datain[111:108] ^ 12);
  assign w101[51] = |(datain[107:104] ^ 13);
  assign w101[52] = |(datain[103:100] ^ 2);
  assign w101[53] = |(datain[99:96] ^ 1);
  assign w101[54] = |(datain[95:92] ^ 7);
  assign w101[55] = |(datain[91:88] ^ 2);
  assign w101[56] = |(datain[87:84] ^ 0);
  assign w101[57] = |(datain[83:80] ^ 10);
  assign w101[58] = |(datain[79:76] ^ 9);
  assign w101[59] = |(datain[75:72] ^ 0);
  assign w101[60] = |(datain[71:68] ^ 9);
  assign w101[61] = |(datain[67:64] ^ 0);
  assign w101[62] = |(datain[63:60] ^ 9);
  assign w101[63] = |(datain[59:56] ^ 0);
  assign w101[64] = |(datain[55:52] ^ 11);
  assign w101[65] = |(datain[51:48] ^ 8);
  assign w101[66] = |(datain[47:44] ^ 0);
  assign w101[67] = |(datain[43:40] ^ 1);
  assign w101[68] = |(datain[39:36] ^ 5);
  assign w101[69] = |(datain[35:32] ^ 7);
  assign w101[70] = |(datain[31:28] ^ 11);
  assign w101[71] = |(datain[27:24] ^ 1);
  assign w101[72] = |(datain[23:20] ^ 1);
  assign w101[73] = |(datain[19:16] ^ 13);
  assign comp[101] = ~(|w101);
  wire [74-1:0] w102;
  assign w102[0] = |(datain[311:308] ^ 11);
  assign w102[1] = |(datain[307:304] ^ 8);
  assign w102[2] = |(datain[303:300] ^ 0);
  assign w102[3] = |(datain[299:296] ^ 0);
  assign w102[4] = |(datain[295:292] ^ 4);
  assign w102[5] = |(datain[291:288] ^ 2);
  assign w102[6] = |(datain[287:284] ^ 14);
  assign w102[7] = |(datain[283:280] ^ 8);
  assign w102[8] = |(datain[279:276] ^ 2);
  assign w102[9] = |(datain[275:272] ^ 11);
  assign w102[10] = |(datain[271:268] ^ 0);
  assign w102[11] = |(datain[267:264] ^ 0);
  assign w102[12] = |(datain[263:260] ^ 8);
  assign w102[13] = |(datain[259:256] ^ 13);
  assign w102[14] = |(datain[255:252] ^ 9);
  assign w102[15] = |(datain[251:248] ^ 6);
  assign w102[16] = |(datain[247:244] ^ 15);
  assign w102[17] = |(datain[243:240] ^ 14);
  assign w102[18] = |(datain[239:236] ^ 0);
  assign w102[19] = |(datain[235:232] ^ 1);
  assign w102[20] = |(datain[231:228] ^ 11);
  assign w102[21] = |(datain[227:224] ^ 9);
  assign w102[22] = |(datain[223:220] ^ 0);
  assign w102[23] = |(datain[219:216] ^ 5);
  assign w102[24] = |(datain[215:212] ^ 0);
  assign w102[25] = |(datain[211:208] ^ 0);
  assign w102[26] = |(datain[207:204] ^ 11);
  assign w102[27] = |(datain[203:200] ^ 4);
  assign w102[28] = |(datain[199:196] ^ 4);
  assign w102[29] = |(datain[195:192] ^ 0);
  assign w102[30] = |(datain[191:188] ^ 12);
  assign w102[31] = |(datain[187:184] ^ 13);
  assign w102[32] = |(datain[183:180] ^ 2);
  assign w102[33] = |(datain[179:176] ^ 1);
  assign w102[34] = |(datain[175:172] ^ 15);
  assign w102[35] = |(datain[171:168] ^ 14);
  assign w102[36] = |(datain[167:164] ^ 8);
  assign w102[37] = |(datain[163:160] ^ 6);
  assign w102[38] = |(datain[159:156] ^ 0);
  assign w102[39] = |(datain[155:152] ^ 5);
  assign w102[40] = |(datain[151:148] ^ 0);
  assign w102[41] = |(datain[147:144] ^ 2);
  assign w102[42] = |(datain[143:140] ^ 5);
  assign w102[43] = |(datain[139:136] ^ 10);
  assign w102[44] = |(datain[135:132] ^ 5);
  assign w102[45] = |(datain[131:128] ^ 9);
  assign w102[46] = |(datain[127:124] ^ 11);
  assign w102[47] = |(datain[123:120] ^ 8);
  assign w102[48] = |(datain[119:116] ^ 0);
  assign w102[49] = |(datain[115:112] ^ 1);
  assign w102[50] = |(datain[111:108] ^ 5);
  assign w102[51] = |(datain[107:104] ^ 7);
  assign w102[52] = |(datain[103:100] ^ 12);
  assign w102[53] = |(datain[99:96] ^ 13);
  assign w102[54] = |(datain[95:92] ^ 2);
  assign w102[55] = |(datain[91:88] ^ 1);
  assign w102[56] = |(datain[87:84] ^ 11);
  assign w102[57] = |(datain[83:80] ^ 4);
  assign w102[58] = |(datain[79:76] ^ 3);
  assign w102[59] = |(datain[75:72] ^ 14);
  assign w102[60] = |(datain[71:68] ^ 12);
  assign w102[61] = |(datain[67:64] ^ 13);
  assign w102[62] = |(datain[63:60] ^ 2);
  assign w102[63] = |(datain[59:56] ^ 1);
  assign w102[64] = |(datain[55:52] ^ 8);
  assign w102[65] = |(datain[51:48] ^ 0);
  assign w102[66] = |(datain[47:44] ^ 11);
  assign w102[67] = |(datain[43:40] ^ 14);
  assign w102[68] = |(datain[39:36] ^ 0);
  assign w102[69] = |(datain[35:32] ^ 5);
  assign w102[70] = |(datain[31:28] ^ 0);
  assign w102[71] = |(datain[27:24] ^ 2);
  assign w102[72] = |(datain[23:20] ^ 0);
  assign w102[73] = |(datain[19:16] ^ 1);
  assign comp[102] = ~(|w102);
  wire [74-1:0] w103;
  assign w103[0] = |(datain[311:308] ^ 0);
  assign w103[1] = |(datain[307:304] ^ 2);
  assign w103[2] = |(datain[303:300] ^ 0);
  assign w103[3] = |(datain[299:296] ^ 5);
  assign w103[4] = |(datain[295:292] ^ 0);
  assign w103[5] = |(datain[291:288] ^ 2);
  assign w103[6] = |(datain[287:284] ^ 0);
  assign w103[7] = |(datain[283:280] ^ 0);
  assign w103[8] = |(datain[279:276] ^ 8);
  assign w103[9] = |(datain[275:272] ^ 9);
  assign w103[10] = |(datain[271:268] ^ 0);
  assign w103[11] = |(datain[267:264] ^ 4);
  assign w103[12] = |(datain[263:260] ^ 8);
  assign w103[13] = |(datain[259:256] ^ 13);
  assign w103[14] = |(datain[255:252] ^ 9);
  assign w103[15] = |(datain[251:248] ^ 6);
  assign w103[16] = |(datain[247:244] ^ 15);
  assign w103[17] = |(datain[243:240] ^ 9);
  assign w103[18] = |(datain[239:236] ^ 0);
  assign w103[19] = |(datain[235:232] ^ 1);
  assign w103[20] = |(datain[231:228] ^ 11);
  assign w103[21] = |(datain[227:224] ^ 9);
  assign w103[22] = |(datain[223:220] ^ 0);
  assign w103[23] = |(datain[219:216] ^ 5);
  assign w103[24] = |(datain[215:212] ^ 0);
  assign w103[25] = |(datain[211:208] ^ 0);
  assign w103[26] = |(datain[207:204] ^ 11);
  assign w103[27] = |(datain[203:200] ^ 4);
  assign w103[28] = |(datain[199:196] ^ 4);
  assign w103[29] = |(datain[195:192] ^ 0);
  assign w103[30] = |(datain[191:188] ^ 12);
  assign w103[31] = |(datain[187:184] ^ 13);
  assign w103[32] = |(datain[183:180] ^ 2);
  assign w103[33] = |(datain[179:176] ^ 1);
  assign w103[34] = |(datain[175:172] ^ 5);
  assign w103[35] = |(datain[171:168] ^ 3);
  assign w103[36] = |(datain[167:164] ^ 5);
  assign w103[37] = |(datain[163:160] ^ 5);
  assign w103[38] = |(datain[159:156] ^ 8);
  assign w103[39] = |(datain[155:152] ^ 11);
  assign w103[40] = |(datain[151:148] ^ 1);
  assign w103[41] = |(datain[147:144] ^ 4);
  assign w103[42] = |(datain[143:140] ^ 8);
  assign w103[43] = |(datain[139:136] ^ 1);
  assign w103[44] = |(datain[135:132] ^ 12);
  assign w103[45] = |(datain[131:128] ^ 2);
  assign w103[46] = |(datain[127:124] ^ 0);
  assign w103[47] = |(datain[123:120] ^ 3);
  assign w103[48] = |(datain[119:116] ^ 0);
  assign w103[49] = |(datain[115:112] ^ 1);
  assign w103[50] = |(datain[111:108] ^ 11);
  assign w103[51] = |(datain[107:104] ^ 9);
  assign w103[52] = |(datain[103:100] ^ 1);
  assign w103[53] = |(datain[99:96] ^ 8);
  assign w103[54] = |(datain[95:92] ^ 0);
  assign w103[55] = |(datain[91:88] ^ 5);
  assign w103[56] = |(datain[87:84] ^ 8);
  assign w103[57] = |(datain[83:80] ^ 13);
  assign w103[58] = |(datain[79:76] ^ 11);
  assign w103[59] = |(datain[75:72] ^ 14);
  assign w103[60] = |(datain[71:68] ^ 10);
  assign w103[61] = |(datain[67:64] ^ 0);
  assign w103[62] = |(datain[63:60] ^ 0);
  assign w103[63] = |(datain[59:56] ^ 6);
  assign w103[64] = |(datain[55:52] ^ 8);
  assign w103[65] = |(datain[51:48] ^ 13);
  assign w103[66] = |(datain[47:44] ^ 11);
  assign w103[67] = |(datain[43:40] ^ 6);
  assign w103[68] = |(datain[39:36] ^ 0);
  assign w103[69] = |(datain[35:32] ^ 8);
  assign w103[70] = |(datain[31:28] ^ 0);
  assign w103[71] = |(datain[27:24] ^ 1);
  assign w103[72] = |(datain[23:20] ^ 14);
  assign w103[73] = |(datain[19:16] ^ 8);
  assign comp[103] = ~(|w103);
  wire [74-1:0] w104;
  assign w104[0] = |(datain[311:308] ^ 12);
  assign w104[1] = |(datain[307:304] ^ 13);
  assign w104[2] = |(datain[303:300] ^ 2);
  assign w104[3] = |(datain[299:296] ^ 1);
  assign w104[4] = |(datain[295:292] ^ 12);
  assign w104[5] = |(datain[291:288] ^ 3);
  assign w104[6] = |(datain[287:284] ^ 11);
  assign w104[7] = |(datain[283:280] ^ 4);
  assign w104[8] = |(datain[279:276] ^ 3);
  assign w104[9] = |(datain[275:272] ^ 14);
  assign w104[10] = |(datain[271:268] ^ 12);
  assign w104[11] = |(datain[267:264] ^ 13);
  assign w104[12] = |(datain[263:260] ^ 2);
  assign w104[13] = |(datain[259:256] ^ 1);
  assign w104[14] = |(datain[255:252] ^ 12);
  assign w104[15] = |(datain[251:248] ^ 3);
  assign w104[16] = |(datain[247:244] ^ 11);
  assign w104[17] = |(datain[243:240] ^ 4);
  assign w104[18] = |(datain[239:236] ^ 3);
  assign w104[19] = |(datain[235:232] ^ 15);
  assign w104[20] = |(datain[231:228] ^ 12);
  assign w104[21] = |(datain[227:224] ^ 13);
  assign w104[22] = |(datain[223:220] ^ 2);
  assign w104[23] = |(datain[219:216] ^ 1);
  assign w104[24] = |(datain[215:212] ^ 12);
  assign w104[25] = |(datain[211:208] ^ 3);
  assign w104[26] = |(datain[207:204] ^ 11);
  assign w104[27] = |(datain[203:200] ^ 4);
  assign w104[28] = |(datain[199:196] ^ 4);
  assign w104[29] = |(datain[195:192] ^ 0);
  assign w104[30] = |(datain[191:188] ^ 12);
  assign w104[31] = |(datain[187:184] ^ 13);
  assign w104[32] = |(datain[183:180] ^ 2);
  assign w104[33] = |(datain[179:176] ^ 1);
  assign w104[34] = |(datain[175:172] ^ 12);
  assign w104[35] = |(datain[171:168] ^ 3);
  assign w104[36] = |(datain[167:164] ^ 11);
  assign w104[37] = |(datain[163:160] ^ 8);
  assign w104[38] = |(datain[159:156] ^ 0);
  assign w104[39] = |(datain[155:152] ^ 0);
  assign w104[40] = |(datain[151:148] ^ 4);
  assign w104[41] = |(datain[147:144] ^ 2);
  assign w104[42] = |(datain[143:140] ^ 3);
  assign w104[43] = |(datain[139:136] ^ 3);
  assign w104[44] = |(datain[135:132] ^ 12);
  assign w104[45] = |(datain[131:128] ^ 9);
  assign w104[46] = |(datain[127:124] ^ 3);
  assign w104[47] = |(datain[123:120] ^ 3);
  assign w104[48] = |(datain[119:116] ^ 13);
  assign w104[49] = |(datain[115:112] ^ 2);
  assign w104[50] = |(datain[111:108] ^ 12);
  assign w104[51] = |(datain[107:104] ^ 13);
  assign w104[52] = |(datain[103:100] ^ 2);
  assign w104[53] = |(datain[99:96] ^ 1);
  assign w104[54] = |(datain[95:92] ^ 12);
  assign w104[55] = |(datain[91:88] ^ 3);
  assign w104[56] = |(datain[87:84] ^ 11);
  assign w104[57] = |(datain[83:80] ^ 8);
  assign w104[58] = |(datain[79:76] ^ 0);
  assign w104[59] = |(datain[75:72] ^ 2);
  assign w104[60] = |(datain[71:68] ^ 4);
  assign w104[61] = |(datain[67:64] ^ 2);
  assign w104[62] = |(datain[63:60] ^ 3);
  assign w104[63] = |(datain[59:56] ^ 3);
  assign w104[64] = |(datain[55:52] ^ 12);
  assign w104[65] = |(datain[51:48] ^ 9);
  assign w104[66] = |(datain[47:44] ^ 3);
  assign w104[67] = |(datain[43:40] ^ 3);
  assign w104[68] = |(datain[39:36] ^ 13);
  assign w104[69] = |(datain[35:32] ^ 2);
  assign w104[70] = |(datain[31:28] ^ 12);
  assign w104[71] = |(datain[27:24] ^ 13);
  assign w104[72] = |(datain[23:20] ^ 2);
  assign w104[73] = |(datain[19:16] ^ 1);
  assign comp[104] = ~(|w104);
  wire [76-1:0] w105;
  assign w105[0] = |(datain[311:308] ^ 3);
  assign w105[1] = |(datain[307:304] ^ 13);
  assign w105[2] = |(datain[303:300] ^ 11);
  assign w105[3] = |(datain[299:296] ^ 10);
  assign w105[4] = |(datain[295:292] ^ 1);
  assign w105[5] = |(datain[291:288] ^ 14);
  assign w105[6] = |(datain[287:284] ^ 0);
  assign w105[7] = |(datain[283:280] ^ 5);
  assign w105[8] = |(datain[279:276] ^ 12);
  assign w105[9] = |(datain[275:272] ^ 13);
  assign w105[10] = |(datain[271:268] ^ 2);
  assign w105[11] = |(datain[267:264] ^ 1);
  assign w105[12] = |(datain[263:260] ^ 8);
  assign w105[13] = |(datain[259:256] ^ 11);
  assign w105[14] = |(datain[255:252] ^ 13);
  assign w105[15] = |(datain[251:248] ^ 8);
  assign w105[16] = |(datain[247:244] ^ 11);
  assign w105[17] = |(datain[243:240] ^ 4);
  assign w105[18] = |(datain[239:236] ^ 4);
  assign w105[19] = |(datain[235:232] ^ 0);
  assign w105[20] = |(datain[231:228] ^ 11);
  assign w105[21] = |(datain[227:224] ^ 10);
  assign w105[22] = |(datain[223:220] ^ 0);
  assign w105[23] = |(datain[219:216] ^ 0);
  assign w105[24] = |(datain[215:212] ^ 0);
  assign w105[25] = |(datain[211:208] ^ 1);
  assign w105[26] = |(datain[207:204] ^ 11);
  assign w105[27] = |(datain[203:200] ^ 9);
  assign w105[28] = |(datain[199:196] ^ 0);
  assign w105[29] = |(datain[195:192] ^ 9);
  assign w105[30] = |(datain[191:188] ^ 0);
  assign w105[31] = |(datain[187:184] ^ 2);
  assign w105[32] = |(datain[183:180] ^ 12);
  assign w105[33] = |(datain[179:176] ^ 13);
  assign w105[34] = |(datain[175:172] ^ 2);
  assign w105[35] = |(datain[171:168] ^ 1);
  assign w105[36] = |(datain[167:164] ^ 11);
  assign w105[37] = |(datain[163:160] ^ 4);
  assign w105[38] = |(datain[159:156] ^ 3);
  assign w105[39] = |(datain[155:152] ^ 14);
  assign w105[40] = |(datain[151:148] ^ 12);
  assign w105[41] = |(datain[147:144] ^ 13);
  assign w105[42] = |(datain[143:140] ^ 2);
  assign w105[43] = |(datain[139:136] ^ 1);
  assign w105[44] = |(datain[135:132] ^ 11);
  assign w105[45] = |(datain[131:128] ^ 4);
  assign w105[46] = |(datain[127:124] ^ 2);
  assign w105[47] = |(datain[123:120] ^ 11);
  assign w105[48] = |(datain[119:116] ^ 11);
  assign w105[49] = |(datain[115:112] ^ 9);
  assign w105[50] = |(datain[111:108] ^ 4);
  assign w105[51] = |(datain[107:104] ^ 3);
  assign w105[52] = |(datain[103:100] ^ 5);
  assign w105[53] = |(datain[99:96] ^ 6);
  assign w105[54] = |(datain[95:92] ^ 11);
  assign w105[55] = |(datain[91:88] ^ 10);
  assign w105[56] = |(datain[87:84] ^ 4);
  assign w105[57] = |(datain[83:80] ^ 13);
  assign w105[58] = |(datain[79:76] ^ 4);
  assign w105[59] = |(datain[75:72] ^ 15);
  assign w105[60] = |(datain[71:68] ^ 12);
  assign w105[61] = |(datain[67:64] ^ 13);
  assign w105[62] = |(datain[63:60] ^ 2);
  assign w105[63] = |(datain[59:56] ^ 1);
  assign w105[64] = |(datain[55:52] ^ 3);
  assign w105[65] = |(datain[51:48] ^ 12);
  assign w105[66] = |(datain[47:44] ^ 0);
  assign w105[67] = |(datain[43:40] ^ 0);
  assign w105[68] = |(datain[39:36] ^ 11);
  assign w105[69] = |(datain[35:32] ^ 10);
  assign w105[70] = |(datain[31:28] ^ 12);
  assign w105[71] = |(datain[27:24] ^ 12);
  assign w105[72] = |(datain[23:20] ^ 0);
  assign w105[73] = |(datain[19:16] ^ 2);
  assign w105[74] = |(datain[15:12] ^ 7);
  assign w105[75] = |(datain[11:8] ^ 5);
  assign comp[105] = ~(|w105);
  wire [74-1:0] w106;
  assign w106[0] = |(datain[311:308] ^ 10);
  assign w106[1] = |(datain[307:304] ^ 3);
  assign w106[2] = |(datain[303:300] ^ 9);
  assign w106[3] = |(datain[299:296] ^ 10);
  assign w106[4] = |(datain[295:292] ^ 0);
  assign w106[5] = |(datain[291:288] ^ 3);
  assign w106[6] = |(datain[287:284] ^ 11);
  assign w106[7] = |(datain[283:280] ^ 8);
  assign w106[8] = |(datain[279:276] ^ 0);
  assign w106[9] = |(datain[275:272] ^ 0);
  assign w106[10] = |(datain[271:268] ^ 4);
  assign w106[11] = |(datain[267:264] ^ 2);
  assign w106[12] = |(datain[263:260] ^ 3);
  assign w106[13] = |(datain[259:256] ^ 3);
  assign w106[14] = |(datain[255:252] ^ 12);
  assign w106[15] = |(datain[251:248] ^ 9);
  assign w106[16] = |(datain[247:244] ^ 9);
  assign w106[17] = |(datain[243:240] ^ 9);
  assign w106[18] = |(datain[239:236] ^ 12);
  assign w106[19] = |(datain[235:232] ^ 13);
  assign w106[20] = |(datain[231:228] ^ 2);
  assign w106[21] = |(datain[227:224] ^ 1);
  assign w106[22] = |(datain[223:220] ^ 11);
  assign w106[23] = |(datain[219:216] ^ 4);
  assign w106[24] = |(datain[215:212] ^ 4);
  assign w106[25] = |(datain[211:208] ^ 0);
  assign w106[26] = |(datain[207:204] ^ 5);
  assign w106[27] = |(datain[203:200] ^ 10);
  assign w106[28] = |(datain[199:196] ^ 5);
  assign w106[29] = |(datain[195:192] ^ 9);
  assign w106[30] = |(datain[191:188] ^ 12);
  assign w106[31] = |(datain[187:184] ^ 13);
  assign w106[32] = |(datain[183:180] ^ 2);
  assign w106[33] = |(datain[179:176] ^ 1);
  assign w106[34] = |(datain[175:172] ^ 5);
  assign w106[35] = |(datain[171:168] ^ 10);
  assign w106[36] = |(datain[167:164] ^ 5);
  assign w106[37] = |(datain[163:160] ^ 9);
  assign w106[38] = |(datain[159:156] ^ 8);
  assign w106[39] = |(datain[155:152] ^ 0);
  assign w106[40] = |(datain[151:148] ^ 12);
  assign w106[41] = |(datain[147:144] ^ 6);
  assign w106[42] = |(datain[143:140] ^ 12);
  assign w106[43] = |(datain[139:136] ^ 8);
  assign w106[44] = |(datain[135:132] ^ 11);
  assign w106[45] = |(datain[131:128] ^ 8);
  assign w106[46] = |(datain[127:124] ^ 0);
  assign w106[47] = |(datain[123:120] ^ 1);
  assign w106[48] = |(datain[119:116] ^ 5);
  assign w106[49] = |(datain[115:112] ^ 7);
  assign w106[50] = |(datain[111:108] ^ 12);
  assign w106[51] = |(datain[107:104] ^ 13);
  assign w106[52] = |(datain[103:100] ^ 2);
  assign w106[53] = |(datain[99:96] ^ 1);
  assign w106[54] = |(datain[95:92] ^ 11);
  assign w106[55] = |(datain[91:88] ^ 4);
  assign w106[56] = |(datain[87:84] ^ 3);
  assign w106[57] = |(datain[83:80] ^ 14);
  assign w106[58] = |(datain[79:76] ^ 12);
  assign w106[59] = |(datain[75:72] ^ 13);
  assign w106[60] = |(datain[71:68] ^ 2);
  assign w106[61] = |(datain[67:64] ^ 1);
  assign w106[62] = |(datain[63:60] ^ 0);
  assign w106[63] = |(datain[59:56] ^ 7);
  assign w106[64] = |(datain[55:52] ^ 1);
  assign w106[65] = |(datain[51:48] ^ 15);
  assign w106[66] = |(datain[47:44] ^ 5);
  assign w106[67] = |(datain[43:40] ^ 14);
  assign w106[68] = |(datain[39:36] ^ 5);
  assign w106[69] = |(datain[35:32] ^ 15);
  assign w106[70] = |(datain[31:28] ^ 5);
  assign w106[71] = |(datain[27:24] ^ 10);
  assign w106[72] = |(datain[23:20] ^ 5);
  assign w106[73] = |(datain[19:16] ^ 9);
  assign comp[106] = ~(|w106);
  wire [74-1:0] w107;
  assign w107[0] = |(datain[311:308] ^ 1);
  assign w107[1] = |(datain[307:304] ^ 0);
  assign w107[2] = |(datain[303:300] ^ 11);
  assign w107[3] = |(datain[299:296] ^ 8);
  assign w107[4] = |(datain[295:292] ^ 0);
  assign w107[5] = |(datain[291:288] ^ 0);
  assign w107[6] = |(datain[287:284] ^ 4);
  assign w107[7] = |(datain[283:280] ^ 2);
  assign w107[8] = |(datain[279:276] ^ 8);
  assign w107[9] = |(datain[275:272] ^ 11);
  assign w107[10] = |(datain[271:268] ^ 12);
  assign w107[11] = |(datain[267:264] ^ 10);
  assign w107[12] = |(datain[263:260] ^ 12);
  assign w107[13] = |(datain[259:256] ^ 13);
  assign w107[14] = |(datain[255:252] ^ 2);
  assign w107[15] = |(datain[251:248] ^ 1);
  assign w107[16] = |(datain[247:244] ^ 11);
  assign w107[17] = |(datain[243:240] ^ 4);
  assign w107[18] = |(datain[239:236] ^ 4);
  assign w107[19] = |(datain[235:232] ^ 0);
  assign w107[20] = |(datain[231:228] ^ 8);
  assign w107[21] = |(datain[227:224] ^ 11);
  assign w107[22] = |(datain[223:220] ^ 13);
  assign w107[23] = |(datain[219:216] ^ 7);
  assign w107[24] = |(datain[215:212] ^ 11);
  assign w107[25] = |(datain[211:208] ^ 9);
  assign w107[26] = |(datain[207:204] ^ 1);
  assign w107[27] = |(datain[203:200] ^ 8);
  assign w107[28] = |(datain[199:196] ^ 0);
  assign w107[29] = |(datain[195:192] ^ 0);
  assign w107[30] = |(datain[191:188] ^ 12);
  assign w107[31] = |(datain[187:184] ^ 13);
  assign w107[32] = |(datain[183:180] ^ 2);
  assign w107[33] = |(datain[179:176] ^ 1);
  assign w107[34] = |(datain[175:172] ^ 5);
  assign w107[35] = |(datain[171:168] ^ 10);
  assign w107[36] = |(datain[167:164] ^ 5);
  assign w107[37] = |(datain[163:160] ^ 9);
  assign w107[38] = |(datain[159:156] ^ 5);
  assign w107[39] = |(datain[155:152] ^ 8);
  assign w107[40] = |(datain[151:148] ^ 4);
  assign w107[41] = |(datain[147:144] ^ 0);
  assign w107[42] = |(datain[143:140] ^ 12);
  assign w107[43] = |(datain[139:136] ^ 13);
  assign w107[44] = |(datain[135:132] ^ 2);
  assign w107[45] = |(datain[131:128] ^ 1);
  assign w107[46] = |(datain[127:124] ^ 11);
  assign w107[47] = |(datain[123:120] ^ 4);
  assign w107[48] = |(datain[119:116] ^ 3);
  assign w107[49] = |(datain[115:112] ^ 14);
  assign w107[50] = |(datain[111:108] ^ 12);
  assign w107[51] = |(datain[107:104] ^ 13);
  assign w107[52] = |(datain[103:100] ^ 2);
  assign w107[53] = |(datain[99:96] ^ 1);
  assign w107[54] = |(datain[95:92] ^ 5);
  assign w107[55] = |(datain[91:88] ^ 10);
  assign w107[56] = |(datain[87:84] ^ 1);
  assign w107[57] = |(datain[83:80] ^ 15);
  assign w107[58] = |(datain[79:76] ^ 5);
  assign w107[59] = |(datain[75:72] ^ 9);
  assign w107[60] = |(datain[71:68] ^ 5);
  assign w107[61] = |(datain[67:64] ^ 8);
  assign w107[62] = |(datain[63:60] ^ 12);
  assign w107[63] = |(datain[59:56] ^ 13);
  assign w107[64] = |(datain[55:52] ^ 2);
  assign w107[65] = |(datain[51:48] ^ 1);
  assign w107[66] = |(datain[47:44] ^ 5);
  assign w107[67] = |(datain[43:40] ^ 8);
  assign w107[68] = |(datain[39:36] ^ 5);
  assign w107[69] = |(datain[35:32] ^ 10);
  assign w107[70] = |(datain[31:28] ^ 1);
  assign w107[71] = |(datain[27:24] ^ 15);
  assign w107[72] = |(datain[23:20] ^ 12);
  assign w107[73] = |(datain[19:16] ^ 13);
  assign comp[107] = ~(|w107);
  wire [76-1:0] w108;
  assign w108[0] = |(datain[311:308] ^ 0);
  assign w108[1] = |(datain[307:304] ^ 2);
  assign w108[2] = |(datain[303:300] ^ 3);
  assign w108[3] = |(datain[299:296] ^ 13);
  assign w108[4] = |(datain[295:292] ^ 11);
  assign w108[5] = |(datain[291:288] ^ 10);
  assign w108[6] = |(datain[287:284] ^ 9);
  assign w108[7] = |(datain[283:280] ^ 14);
  assign w108[8] = |(datain[279:276] ^ 0);
  assign w108[9] = |(datain[275:272] ^ 0);
  assign w108[10] = |(datain[271:268] ^ 12);
  assign w108[11] = |(datain[267:264] ^ 13);
  assign w108[12] = |(datain[263:260] ^ 2);
  assign w108[13] = |(datain[259:256] ^ 1);
  assign w108[14] = |(datain[255:252] ^ 9);
  assign w108[15] = |(datain[251:248] ^ 3);
  assign w108[16] = |(datain[247:244] ^ 11);
  assign w108[17] = |(datain[243:240] ^ 4);
  assign w108[18] = |(datain[239:236] ^ 4);
  assign w108[19] = |(datain[235:232] ^ 0);
  assign w108[20] = |(datain[231:228] ^ 11);
  assign w108[21] = |(datain[227:224] ^ 10);
  assign w108[22] = |(datain[223:220] ^ 0);
  assign w108[23] = |(datain[219:216] ^ 0);
  assign w108[24] = |(datain[215:212] ^ 0);
  assign w108[25] = |(datain[211:208] ^ 1);
  assign w108[26] = |(datain[207:204] ^ 11);
  assign w108[27] = |(datain[203:200] ^ 9);
  assign w108[28] = |(datain[199:196] ^ 7);
  assign w108[29] = |(datain[195:192] ^ 15);
  assign w108[30] = |(datain[191:188] ^ 0);
  assign w108[31] = |(datain[187:184] ^ 2);
  assign w108[32] = |(datain[183:180] ^ 12);
  assign w108[33] = |(datain[179:176] ^ 13);
  assign w108[34] = |(datain[175:172] ^ 2);
  assign w108[35] = |(datain[171:168] ^ 1);
  assign w108[36] = |(datain[167:164] ^ 11);
  assign w108[37] = |(datain[163:160] ^ 4);
  assign w108[38] = |(datain[159:156] ^ 3);
  assign w108[39] = |(datain[155:152] ^ 14);
  assign w108[40] = |(datain[151:148] ^ 12);
  assign w108[41] = |(datain[147:144] ^ 13);
  assign w108[42] = |(datain[143:140] ^ 2);
  assign w108[43] = |(datain[139:136] ^ 1);
  assign w108[44] = |(datain[135:132] ^ 11);
  assign w108[45] = |(datain[131:128] ^ 4);
  assign w108[46] = |(datain[127:124] ^ 4);
  assign w108[47] = |(datain[123:120] ^ 15);
  assign w108[48] = |(datain[119:116] ^ 14);
  assign w108[49] = |(datain[115:112] ^ 11);
  assign w108[50] = |(datain[111:108] ^ 13);
  assign w108[51] = |(datain[107:104] ^ 10);
  assign w108[52] = |(datain[103:100] ^ 11);
  assign w108[53] = |(datain[99:96] ^ 10);
  assign w108[54] = |(datain[95:92] ^ 5);
  assign w108[55] = |(datain[91:88] ^ 8);
  assign w108[56] = |(datain[87:84] ^ 0);
  assign w108[57] = |(datain[83:80] ^ 2);
  assign w108[58] = |(datain[79:76] ^ 11);
  assign w108[59] = |(datain[75:72] ^ 4);
  assign w108[60] = |(datain[71:68] ^ 0);
  assign w108[61] = |(datain[67:64] ^ 9);
  assign w108[62] = |(datain[63:60] ^ 15);
  assign w108[63] = |(datain[59:56] ^ 14);
  assign w108[64] = |(datain[55:52] ^ 12);
  assign w108[65] = |(datain[51:48] ^ 6);
  assign w108[66] = |(datain[47:44] ^ 12);
  assign w108[67] = |(datain[43:40] ^ 13);
  assign w108[68] = |(datain[39:36] ^ 2);
  assign w108[69] = |(datain[35:32] ^ 1);
  assign w108[70] = |(datain[31:28] ^ 12);
  assign w108[71] = |(datain[27:24] ^ 13);
  assign w108[72] = |(datain[23:20] ^ 2);
  assign w108[73] = |(datain[19:16] ^ 0);
  assign w108[74] = |(datain[15:12] ^ 2);
  assign w108[75] = |(datain[11:8] ^ 10);
  assign comp[108] = ~(|w108);
  wire [76-1:0] w109;
  assign w109[0] = |(datain[311:308] ^ 8);
  assign w109[1] = |(datain[307:304] ^ 11);
  assign w109[2] = |(datain[303:300] ^ 0);
  assign w109[3] = |(datain[299:296] ^ 4);
  assign w109[4] = |(datain[295:292] ^ 8);
  assign w109[5] = |(datain[291:288] ^ 13);
  assign w109[6] = |(datain[287:284] ^ 11);
  assign w109[7] = |(datain[283:280] ^ 14);
  assign w109[8] = |(datain[279:276] ^ 0);
  assign w109[9] = |(datain[275:272] ^ 14);
  assign w109[10] = |(datain[271:268] ^ 0);
  assign w109[11] = |(datain[267:264] ^ 1);
  assign w109[12] = |(datain[263:260] ^ 0);
  assign w109[13] = |(datain[259:256] ^ 3);
  assign w109[14] = |(datain[255:252] ^ 0);
  assign w109[15] = |(datain[251:248] ^ 5);
  assign w109[16] = |(datain[247:244] ^ 5);
  assign w109[17] = |(datain[243:240] ^ 0);
  assign w109[18] = |(datain[239:236] ^ 8);
  assign w109[19] = |(datain[235:232] ^ 11);
  assign w109[20] = |(datain[231:228] ^ 13);
  assign w109[21] = |(datain[227:224] ^ 4);
  assign w109[22] = |(datain[223:220] ^ 11);
  assign w109[23] = |(datain[219:216] ^ 4);
  assign w109[24] = |(datain[215:212] ^ 4);
  assign w109[25] = |(datain[211:208] ^ 0);
  assign w109[26] = |(datain[207:204] ^ 11);
  assign w109[27] = |(datain[203:200] ^ 9);
  assign w109[28] = |(datain[199:196] ^ 0);
  assign w109[29] = |(datain[195:192] ^ 2);
  assign w109[30] = |(datain[191:188] ^ 0);
  assign w109[31] = |(datain[187:184] ^ 0);
  assign w109[32] = |(datain[183:180] ^ 12);
  assign w109[33] = |(datain[179:176] ^ 13);
  assign w109[34] = |(datain[175:172] ^ 2);
  assign w109[35] = |(datain[171:168] ^ 1);
  assign w109[36] = |(datain[167:164] ^ 4);
  assign w109[37] = |(datain[163:160] ^ 6);
  assign w109[38] = |(datain[159:156] ^ 4);
  assign w109[39] = |(datain[155:152] ^ 6);
  assign w109[40] = |(datain[151:148] ^ 5);
  assign w109[41] = |(datain[147:144] ^ 8);
  assign w109[42] = |(datain[143:140] ^ 5);
  assign w109[43] = |(datain[139:136] ^ 9);
  assign w109[44] = |(datain[135:132] ^ 14);
  assign w109[45] = |(datain[131:128] ^ 2);
  assign w109[46] = |(datain[127:124] ^ 14);
  assign w109[47] = |(datain[123:120] ^ 7);
  assign w109[48] = |(datain[119:116] ^ 11);
  assign w109[49] = |(datain[115:112] ^ 8);
  assign w109[50] = |(datain[111:108] ^ 0);
  assign w109[51] = |(datain[107:104] ^ 0);
  assign w109[52] = |(datain[103:100] ^ 4);
  assign w109[53] = |(datain[99:96] ^ 2);
  assign w109[54] = |(datain[95:92] ^ 11);
  assign w109[55] = |(datain[91:88] ^ 9);
  assign w109[56] = |(datain[87:84] ^ 0);
  assign w109[57] = |(datain[83:80] ^ 0);
  assign w109[58] = |(datain[79:76] ^ 0);
  assign w109[59] = |(datain[75:72] ^ 0);
  assign w109[60] = |(datain[71:68] ^ 11);
  assign w109[61] = |(datain[67:64] ^ 10);
  assign w109[62] = |(datain[63:60] ^ 0);
  assign w109[63] = |(datain[59:56] ^ 0);
  assign w109[64] = |(datain[55:52] ^ 0);
  assign w109[65] = |(datain[51:48] ^ 0);
  assign w109[66] = |(datain[47:44] ^ 12);
  assign w109[67] = |(datain[43:40] ^ 13);
  assign w109[68] = |(datain[39:36] ^ 2);
  assign w109[69] = |(datain[35:32] ^ 1);
  assign w109[70] = |(datain[31:28] ^ 8);
  assign w109[71] = |(datain[27:24] ^ 13);
  assign w109[72] = |(datain[23:20] ^ 9);
  assign w109[73] = |(datain[19:16] ^ 6);
  assign w109[74] = |(datain[15:12] ^ 3);
  assign w109[75] = |(datain[11:8] ^ 7);
  assign comp[109] = ~(|w109);
  wire [76-1:0] w110;
  assign w110[0] = |(datain[311:308] ^ 10);
  assign w110[1] = |(datain[307:304] ^ 4);
  assign w110[2] = |(datain[303:300] ^ 0);
  assign w110[3] = |(datain[299:296] ^ 8);
  assign w110[4] = |(datain[295:292] ^ 2);
  assign w110[5] = |(datain[291:288] ^ 14);
  assign w110[6] = |(datain[287:284] ^ 8);
  assign w110[7] = |(datain[283:280] ^ 11);
  assign w110[8] = |(datain[279:276] ^ 9);
  assign w110[9] = |(datain[275:272] ^ 6);
  assign w110[10] = |(datain[271:268] ^ 10);
  assign w110[11] = |(datain[267:264] ^ 6);
  assign w110[12] = |(datain[263:260] ^ 0);
  assign w110[13] = |(datain[259:256] ^ 8);
  assign w110[14] = |(datain[255:252] ^ 12);
  assign w110[15] = |(datain[251:248] ^ 13);
  assign w110[16] = |(datain[247:244] ^ 7);
  assign w110[17] = |(datain[243:240] ^ 9);
  assign w110[18] = |(datain[239:236] ^ 14);
  assign w110[19] = |(datain[235:232] ^ 8);
  assign w110[20] = |(datain[231:228] ^ 2);
  assign w110[21] = |(datain[227:224] ^ 0);
  assign w110[22] = |(datain[223:220] ^ 0);
  assign w110[23] = |(datain[219:216] ^ 0);
  assign w110[24] = |(datain[215:212] ^ 12);
  assign w110[25] = |(datain[211:208] ^ 3);
  assign w110[26] = |(datain[207:204] ^ 5);
  assign w110[27] = |(datain[203:200] ^ 0);
  assign w110[28] = |(datain[199:196] ^ 11);
  assign w110[29] = |(datain[195:192] ^ 4);
  assign w110[30] = |(datain[191:188] ^ 4);
  assign w110[31] = |(datain[187:184] ^ 0);
  assign w110[32] = |(datain[183:180] ^ 12);
  assign w110[33] = |(datain[179:176] ^ 13);
  assign w110[34] = |(datain[175:172] ^ 7);
  assign w110[35] = |(datain[171:168] ^ 9);
  assign w110[36] = |(datain[167:164] ^ 3);
  assign w110[37] = |(datain[163:160] ^ 11);
  assign w110[38] = |(datain[159:156] ^ 12);
  assign w110[39] = |(datain[155:152] ^ 1);
  assign w110[40] = |(datain[151:148] ^ 7);
  assign w110[41] = |(datain[147:144] ^ 4);
  assign w110[42] = |(datain[143:140] ^ 0);
  assign w110[43] = |(datain[139:136] ^ 1);
  assign w110[44] = |(datain[135:132] ^ 15);
  assign w110[45] = |(datain[131:128] ^ 9);
  assign w110[46] = |(datain[127:124] ^ 5);
  assign w110[47] = |(datain[123:120] ^ 8);
  assign w110[48] = |(datain[119:116] ^ 12);
  assign w110[49] = |(datain[115:112] ^ 3);
  assign w110[50] = |(datain[111:108] ^ 2);
  assign w110[51] = |(datain[107:104] ^ 14);
  assign w110[52] = |(datain[103:100] ^ 8);
  assign w110[53] = |(datain[99:96] ^ 15);
  assign w110[54] = |(datain[95:92] ^ 8);
  assign w110[55] = |(datain[91:88] ^ 6);
  assign w110[56] = |(datain[87:84] ^ 8);
  assign w110[57] = |(datain[83:80] ^ 12);
  assign w110[58] = |(datain[79:76] ^ 0);
  assign w110[59] = |(datain[75:72] ^ 8);
  assign w110[60] = |(datain[71:68] ^ 5);
  assign w110[61] = |(datain[67:64] ^ 0);
  assign w110[62] = |(datain[63:60] ^ 5);
  assign w110[63] = |(datain[59:56] ^ 3);
  assign w110[64] = |(datain[55:52] ^ 5);
  assign w110[65] = |(datain[51:48] ^ 1);
  assign w110[66] = |(datain[47:44] ^ 5);
  assign w110[67] = |(datain[43:40] ^ 2);
  assign w110[68] = |(datain[39:36] ^ 5);
  assign w110[69] = |(datain[35:32] ^ 7);
  assign w110[70] = |(datain[31:28] ^ 5);
  assign w110[71] = |(datain[27:24] ^ 6);
  assign w110[72] = |(datain[23:20] ^ 1);
  assign w110[73] = |(datain[19:16] ^ 14);
  assign w110[74] = |(datain[15:12] ^ 0);
  assign w110[75] = |(datain[11:8] ^ 6);
  assign comp[110] = ~(|w110);
  wire [76-1:0] w111;
  assign w111[0] = |(datain[311:308] ^ 11);
  assign w111[1] = |(datain[307:304] ^ 9);
  assign w111[2] = |(datain[303:300] ^ 10);
  assign w111[3] = |(datain[299:296] ^ 14);
  assign w111[4] = |(datain[295:292] ^ 0);
  assign w111[5] = |(datain[291:288] ^ 7);
  assign w111[6] = |(datain[287:284] ^ 3);
  assign w111[7] = |(datain[283:280] ^ 0);
  assign w111[8] = |(datain[279:276] ^ 0);
  assign w111[9] = |(datain[275:272] ^ 4);
  assign w111[10] = |(datain[271:268] ^ 4);
  assign w111[11] = |(datain[267:264] ^ 6);
  assign w111[12] = |(datain[263:260] ^ 14);
  assign w111[13] = |(datain[259:256] ^ 2);
  assign w111[14] = |(datain[255:252] ^ 15);
  assign w111[15] = |(datain[251:248] ^ 11);
  assign w111[16] = |(datain[247:244] ^ 11);
  assign w111[17] = |(datain[243:240] ^ 4);
  assign w111[18] = |(datain[239:236] ^ 4);
  assign w111[19] = |(datain[235:232] ^ 0);
  assign w111[20] = |(datain[231:228] ^ 11);
  assign w111[21] = |(datain[227:224] ^ 9);
  assign w111[22] = |(datain[223:220] ^ 10);
  assign w111[23] = |(datain[219:216] ^ 14);
  assign w111[24] = |(datain[215:212] ^ 0);
  assign w111[25] = |(datain[211:208] ^ 7);
  assign w111[26] = |(datain[207:204] ^ 11);
  assign w111[27] = |(datain[203:200] ^ 10);
  assign w111[28] = |(datain[199:196] ^ 13);
  assign w111[29] = |(datain[195:192] ^ 0);
  assign w111[30] = |(datain[191:188] ^ 0);
  assign w111[31] = |(datain[187:184] ^ 7);
  assign w111[32] = |(datain[183:180] ^ 12);
  assign w111[33] = |(datain[179:176] ^ 13);
  assign w111[34] = |(datain[175:172] ^ 2);
  assign w111[35] = |(datain[171:168] ^ 1);
  assign w111[36] = |(datain[167:164] ^ 14);
  assign w111[37] = |(datain[163:160] ^ 8);
  assign w111[38] = |(datain[159:156] ^ 7);
  assign w111[39] = |(datain[155:152] ^ 9);
  assign w111[40] = |(datain[151:148] ^ 0);
  assign w111[41] = |(datain[147:144] ^ 0);
  assign w111[42] = |(datain[143:140] ^ 11);
  assign w111[43] = |(datain[139:136] ^ 15);
  assign w111[44] = |(datain[135:132] ^ 11);
  assign w111[45] = |(datain[131:128] ^ 2);
  assign w111[46] = |(datain[127:124] ^ 0);
  assign w111[47] = |(datain[123:120] ^ 7);
  assign w111[48] = |(datain[119:116] ^ 11);
  assign w111[49] = |(datain[115:112] ^ 9);
  assign w111[50] = |(datain[111:108] ^ 1);
  assign w111[51] = |(datain[107:104] ^ 14);
  assign w111[52] = |(datain[103:100] ^ 0);
  assign w111[53] = |(datain[99:96] ^ 0);
  assign w111[54] = |(datain[95:92] ^ 5);
  assign w111[55] = |(datain[91:88] ^ 1);
  assign w111[56] = |(datain[87:84] ^ 5);
  assign w111[57] = |(datain[83:80] ^ 7);
  assign w111[58] = |(datain[79:76] ^ 11);
  assign w111[59] = |(datain[75:72] ^ 9);
  assign w111[60] = |(datain[71:68] ^ 2);
  assign w111[61] = |(datain[67:64] ^ 8);
  assign w111[62] = |(datain[63:60] ^ 0);
  assign w111[63] = |(datain[59:56] ^ 0);
  assign w111[64] = |(datain[55:52] ^ 14);
  assign w111[65] = |(datain[51:48] ^ 8);
  assign w111[66] = |(datain[47:44] ^ 13);
  assign w111[67] = |(datain[43:40] ^ 10);
  assign w111[68] = |(datain[39:36] ^ 0);
  assign w111[69] = |(datain[35:32] ^ 3);
  assign w111[70] = |(datain[31:28] ^ 11);
  assign w111[71] = |(datain[27:24] ^ 14);
  assign w111[72] = |(datain[23:20] ^ 4);
  assign w111[73] = |(datain[19:16] ^ 4);
  assign w111[74] = |(datain[15:12] ^ 0);
  assign w111[75] = |(datain[11:8] ^ 7);
  assign comp[111] = ~(|w111);
  wire [76-1:0] w112;
  assign w112[0] = |(datain[311:308] ^ 0);
  assign w112[1] = |(datain[307:304] ^ 14);
  assign w112[2] = |(datain[303:300] ^ 0);
  assign w112[3] = |(datain[299:296] ^ 0);
  assign w112[4] = |(datain[295:292] ^ 3);
  assign w112[5] = |(datain[291:288] ^ 12);
  assign w112[6] = |(datain[287:284] ^ 0);
  assign w112[7] = |(datain[283:280] ^ 6);
  assign w112[8] = |(datain[279:276] ^ 7);
  assign w112[9] = |(datain[275:272] ^ 5);
  assign w112[10] = |(datain[271:268] ^ 0);
  assign w112[11] = |(datain[267:264] ^ 8);
  assign w112[12] = |(datain[263:260] ^ 11);
  assign w112[13] = |(datain[259:256] ^ 4);
  assign w112[14] = |(datain[255:252] ^ 0);
  assign w112[15] = |(datain[251:248] ^ 9);
  assign w112[16] = |(datain[247:244] ^ 11);
  assign w112[17] = |(datain[243:240] ^ 10);
  assign w112[18] = |(datain[239:236] ^ 12);
  assign w112[19] = |(datain[235:232] ^ 8);
  assign w112[20] = |(datain[231:228] ^ 0);
  assign w112[21] = |(datain[227:224] ^ 1);
  assign w112[22] = |(datain[223:220] ^ 14);
  assign w112[23] = |(datain[219:216] ^ 8);
  assign w112[24] = |(datain[215:212] ^ 0);
  assign w112[25] = |(datain[211:208] ^ 2);
  assign w112[26] = |(datain[207:204] ^ 0);
  assign w112[27] = |(datain[203:200] ^ 0);
  assign w112[28] = |(datain[199:196] ^ 12);
  assign w112[29] = |(datain[195:192] ^ 13);
  assign w112[30] = |(datain[191:188] ^ 2);
  assign w112[31] = |(datain[187:184] ^ 0);
  assign w112[32] = |(datain[183:180] ^ 12);
  assign w112[33] = |(datain[179:176] ^ 13);
  assign w112[34] = |(datain[175:172] ^ 2);
  assign w112[35] = |(datain[171:168] ^ 1);
  assign w112[36] = |(datain[167:164] ^ 12);
  assign w112[37] = |(datain[163:160] ^ 3);
  assign w112[38] = |(datain[159:156] ^ 0);
  assign w112[39] = |(datain[155:152] ^ 10);
  assign w112[40] = |(datain[151:148] ^ 0);
  assign w112[41] = |(datain[147:144] ^ 13);
  assign w112[42] = |(datain[143:140] ^ 4);
  assign w112[43] = |(datain[139:136] ^ 1);
  assign w112[44] = |(datain[135:132] ^ 6);
  assign w112[45] = |(datain[131:128] ^ 3);
  assign w112[46] = |(datain[127:124] ^ 7);
  assign w112[47] = |(datain[123:120] ^ 5);
  assign w112[48] = |(datain[119:116] ^ 7);
  assign w112[49] = |(datain[115:112] ^ 2);
  assign w112[50] = |(datain[111:108] ^ 6);
  assign w112[51] = |(datain[107:104] ^ 5);
  assign w112[52] = |(datain[103:100] ^ 7);
  assign w112[53] = |(datain[99:96] ^ 6);
  assign w112[54] = |(datain[95:92] ^ 2);
  assign w112[55] = |(datain[91:88] ^ 0);
  assign w112[56] = |(datain[87:84] ^ 7);
  assign w112[57] = |(datain[83:80] ^ 6);
  assign w112[58] = |(datain[79:76] ^ 3);
  assign w112[59] = |(datain[75:72] ^ 1);
  assign w112[60] = |(datain[71:68] ^ 2);
  assign w112[61] = |(datain[67:64] ^ 14);
  assign w112[62] = |(datain[63:60] ^ 3);
  assign w112[63] = |(datain[59:56] ^ 8);
  assign w112[64] = |(datain[55:52] ^ 2);
  assign w112[65] = |(datain[51:48] ^ 0);
  assign w112[66] = |(datain[47:44] ^ 6);
  assign w112[67] = |(datain[43:40] ^ 3);
  assign w112[68] = |(datain[39:36] ^ 6);
  assign w112[69] = |(datain[35:32] ^ 15);
  assign w112[70] = |(datain[31:28] ^ 6);
  assign w112[71] = |(datain[27:24] ^ 4);
  assign w112[72] = |(datain[23:20] ^ 6);
  assign w112[73] = |(datain[19:16] ^ 5);
  assign w112[74] = |(datain[15:12] ^ 6);
  assign w112[75] = |(datain[11:8] ^ 4);
  assign comp[112] = ~(|w112);
  wire [76-1:0] w113;
  assign w113[0] = |(datain[311:308] ^ 10);
  assign w113[1] = |(datain[307:304] ^ 5);
  assign w113[2] = |(datain[303:300] ^ 0);
  assign w113[3] = |(datain[299:296] ^ 1);
  assign w113[4] = |(datain[295:292] ^ 7);
  assign w113[5] = |(datain[291:288] ^ 3);
  assign w113[6] = |(datain[287:284] ^ 0);
  assign w113[7] = |(datain[283:280] ^ 3);
  assign w113[8] = |(datain[279:276] ^ 14);
  assign w113[9] = |(datain[275:272] ^ 9);
  assign w113[10] = |(datain[271:268] ^ 3);
  assign w113[11] = |(datain[267:264] ^ 15);
  assign w113[12] = |(datain[263:260] ^ 0);
  assign w113[13] = |(datain[259:256] ^ 1);
  assign w113[14] = |(datain[255:252] ^ 11);
  assign w113[15] = |(datain[251:248] ^ 9);
  assign w113[16] = |(datain[247:244] ^ 0);
  assign w113[17] = |(datain[243:240] ^ 3);
  assign w113[18] = |(datain[239:236] ^ 0);
  assign w113[19] = |(datain[235:232] ^ 0);
  assign w113[20] = |(datain[231:228] ^ 8);
  assign w113[21] = |(datain[227:224] ^ 13);
  assign w113[22] = |(datain[223:220] ^ 1);
  assign w113[23] = |(datain[219:216] ^ 6);
  assign w113[24] = |(datain[215:212] ^ 4);
  assign w113[25] = |(datain[211:208] ^ 5);
  assign w113[26] = |(datain[207:204] ^ 0);
  assign w113[27] = |(datain[203:200] ^ 1);
  assign w113[28] = |(datain[199:196] ^ 11);
  assign w113[29] = |(datain[195:192] ^ 4);
  assign w113[30] = |(datain[191:188] ^ 4);
  assign w113[31] = |(datain[187:184] ^ 0);
  assign w113[32] = |(datain[183:180] ^ 12);
  assign w113[33] = |(datain[179:176] ^ 13);
  assign w113[34] = |(datain[175:172] ^ 2);
  assign w113[35] = |(datain[171:168] ^ 1);
  assign w113[36] = |(datain[167:164] ^ 14);
  assign w113[37] = |(datain[163:160] ^ 9);
  assign w113[38] = |(datain[159:156] ^ 3);
  assign w113[39] = |(datain[155:152] ^ 1);
  assign w113[40] = |(datain[151:148] ^ 0);
  assign w113[41] = |(datain[147:144] ^ 1);
  assign w113[42] = |(datain[143:140] ^ 0);
  assign w113[43] = |(datain[139:136] ^ 14);
  assign w113[44] = |(datain[135:132] ^ 1);
  assign w113[45] = |(datain[131:128] ^ 15);
  assign w113[46] = |(datain[127:124] ^ 2);
  assign w113[47] = |(datain[123:120] ^ 14);
  assign w113[48] = |(datain[119:116] ^ 8);
  assign w113[49] = |(datain[115:112] ^ 11);
  assign w113[50] = |(datain[111:108] ^ 1);
  assign w113[51] = |(datain[107:104] ^ 14);
  assign w113[52] = |(datain[103:100] ^ 5);
  assign w113[53] = |(datain[99:96] ^ 2);
  assign w113[54] = |(datain[95:92] ^ 0);
  assign w113[55] = |(datain[91:88] ^ 1);
  assign w113[56] = |(datain[87:84] ^ 11);
  assign w113[57] = |(datain[83:80] ^ 8);
  assign w113[58] = |(datain[79:76] ^ 0);
  assign w113[59] = |(datain[75:72] ^ 2);
  assign w113[60] = |(datain[71:68] ^ 4);
  assign w113[61] = |(datain[67:64] ^ 2);
  assign w113[62] = |(datain[63:60] ^ 11);
  assign w113[63] = |(datain[59:56] ^ 9);
  assign w113[64] = |(datain[55:52] ^ 15);
  assign w113[65] = |(datain[51:48] ^ 15);
  assign w113[66] = |(datain[47:44] ^ 15);
  assign w113[67] = |(datain[43:40] ^ 15);
  assign w113[68] = |(datain[39:36] ^ 11);
  assign w113[69] = |(datain[35:32] ^ 10);
  assign w113[70] = |(datain[31:28] ^ 15);
  assign w113[71] = |(datain[27:24] ^ 14);
  assign w113[72] = |(datain[23:20] ^ 15);
  assign w113[73] = |(datain[19:16] ^ 15);
  assign w113[74] = |(datain[15:12] ^ 12);
  assign w113[75] = |(datain[11:8] ^ 13);
  assign comp[113] = ~(|w113);
  wire [32-1:0] w114;
  assign w114[0] = |(datain[311:308] ^ 8);
  assign w114[1] = |(datain[307:304] ^ 12);
  assign w114[2] = |(datain[303:300] ^ 12);
  assign w114[3] = |(datain[299:296] ^ 0);
  assign w114[4] = |(datain[295:292] ^ 4);
  assign w114[5] = |(datain[291:288] ^ 8);
  assign w114[6] = |(datain[287:284] ^ 8);
  assign w114[7] = |(datain[283:280] ^ 14);
  assign w114[8] = |(datain[279:276] ^ 12);
  assign w114[9] = |(datain[275:272] ^ 0);
  assign w114[10] = |(datain[271:268] ^ 2);
  assign w114[11] = |(datain[267:264] ^ 6);
  assign w114[12] = |(datain[263:260] ^ 10);
  assign w114[13] = |(datain[259:256] ^ 1);
  assign w114[14] = |(datain[255:252] ^ 0);
  assign w114[15] = |(datain[251:248] ^ 3);
  assign w114[16] = |(datain[247:244] ^ 0);
  assign w114[17] = |(datain[243:240] ^ 0);
  assign w114[18] = |(datain[239:236] ^ 2);
  assign w114[19] = |(datain[235:232] ^ 13);
  assign w114[20] = |(datain[231:228] ^ 8);
  assign w114[21] = |(datain[227:224] ^ 0);
  assign w114[22] = |(datain[223:220] ^ 0);
  assign w114[23] = |(datain[219:216] ^ 0);
  assign w114[24] = |(datain[215:212] ^ 2);
  assign w114[25] = |(datain[211:208] ^ 6);
  assign w114[26] = |(datain[207:204] ^ 10);
  assign w114[27] = |(datain[203:200] ^ 3);
  assign w114[28] = |(datain[199:196] ^ 0);
  assign w114[29] = |(datain[195:192] ^ 3);
  assign w114[30] = |(datain[191:188] ^ 0);
  assign w114[31] = |(datain[187:184] ^ 0);
  assign comp[114] = ~(|w114);
  wire [28-1:0] w115;
  assign w115[0] = |(datain[311:308] ^ 0);
  assign w115[1] = |(datain[307:304] ^ 4);
  assign w115[2] = |(datain[303:300] ^ 1);
  assign w115[3] = |(datain[299:296] ^ 15);
  assign w115[4] = |(datain[295:292] ^ 3);
  assign w115[5] = |(datain[291:288] ^ 13);
  assign w115[6] = |(datain[287:284] ^ 15);
  assign w115[7] = |(datain[283:280] ^ 0);
  assign w115[8] = |(datain[279:276] ^ 15);
  assign w115[9] = |(datain[275:272] ^ 0);
  assign w115[10] = |(datain[271:268] ^ 7);
  assign w115[11] = |(datain[267:264] ^ 5);
  assign w115[12] = |(datain[263:260] ^ 0);
  assign w115[13] = |(datain[259:256] ^ 5);
  assign w115[14] = |(datain[255:252] ^ 10);
  assign w115[15] = |(datain[251:248] ^ 1);
  assign w115[16] = |(datain[247:244] ^ 0);
  assign w115[17] = |(datain[243:240] ^ 3);
  assign w115[18] = |(datain[239:236] ^ 0);
  assign w115[19] = |(datain[235:232] ^ 1);
  assign w115[20] = |(datain[231:228] ^ 12);
  assign w115[21] = |(datain[227:224] ^ 13);
  assign w115[22] = |(datain[223:220] ^ 0);
  assign w115[23] = |(datain[219:216] ^ 5);
  assign w115[24] = |(datain[215:212] ^ 2);
  assign w115[25] = |(datain[211:208] ^ 6);
  assign w115[26] = |(datain[207:204] ^ 10);
  assign w115[27] = |(datain[203:200] ^ 1);
  assign comp[115] = ~(|w115);
  wire [40-1:0] w116;
  assign w116[0] = |(datain[311:308] ^ 0);
  assign w116[1] = |(datain[307:304] ^ 1);
  assign w116[2] = |(datain[303:300] ^ 2);
  assign w116[3] = |(datain[299:296] ^ 14);
  assign w116[4] = |(datain[295:292] ^ 10);
  assign w116[5] = |(datain[291:288] ^ 3);
  assign w116[6] = |(datain[287:284] ^ 0);
  assign w116[7] = |(datain[283:280] ^ 3);
  assign w116[8] = |(datain[279:276] ^ 0);
  assign w116[9] = |(datain[275:272] ^ 0);
  assign w116[10] = |(datain[271:268] ^ 11);
  assign w116[11] = |(datain[267:264] ^ 4);
  assign w116[12] = |(datain[263:260] ^ 4);
  assign w116[13] = |(datain[259:256] ^ 0);
  assign w116[14] = |(datain[255:252] ^ 0);
  assign w116[15] = |(datain[251:248] ^ 14);
  assign w116[16] = |(datain[247:244] ^ 1);
  assign w116[17] = |(datain[243:240] ^ 15);
  assign w116[18] = |(datain[239:236] ^ 11);
  assign w116[19] = |(datain[235:232] ^ 10);
  assign w116[20] = |(datain[231:228] ^ 0);
  assign w116[21] = |(datain[227:224] ^ 0);
  assign w116[22] = |(datain[223:220] ^ 0);
  assign w116[23] = |(datain[219:216] ^ 4);
  assign w116[24] = |(datain[215:212] ^ 11);
  assign w116[25] = |(datain[211:208] ^ 9);
  assign w116[26] = |(datain[207:204] ^ 0);
  assign w116[27] = |(datain[203:200] ^ 0);
  assign w116[28] = |(datain[199:196] ^ 0);
  assign w116[29] = |(datain[195:192] ^ 4);
  assign w116[30] = |(datain[191:188] ^ 14);
  assign w116[31] = |(datain[187:184] ^ 8);
  assign w116[32] = |(datain[183:180] ^ 14);
  assign w116[33] = |(datain[179:176] ^ 8);
  assign w116[34] = |(datain[175:172] ^ 0);
  assign w116[35] = |(datain[171:168] ^ 0);
  assign w116[36] = |(datain[167:164] ^ 7);
  assign w116[37] = |(datain[163:160] ^ 2);
  assign w116[38] = |(datain[159:156] ^ 3);
  assign w116[39] = |(datain[155:152] ^ 0);
  assign comp[116] = ~(|w116);
  wire [30-1:0] w117;
  assign w117[0] = |(datain[311:308] ^ 11);
  assign w117[1] = |(datain[307:304] ^ 15);
  assign w117[2] = |(datain[303:300] ^ 0);
  assign w117[3] = |(datain[299:296] ^ 0);
  assign w117[4] = |(datain[295:292] ^ 11);
  assign w117[5] = |(datain[291:288] ^ 8);
  assign w117[6] = |(datain[287:284] ^ 2);
  assign w117[7] = |(datain[283:280] ^ 1);
  assign w117[8] = |(datain[279:276] ^ 2);
  assign w117[9] = |(datain[275:272] ^ 5);
  assign w117[10] = |(datain[271:268] ^ 12);
  assign w117[11] = |(datain[267:264] ^ 13);
  assign w117[12] = |(datain[263:260] ^ 2);
  assign w117[13] = |(datain[259:256] ^ 1);
  assign w117[14] = |(datain[255:252] ^ 3);
  assign w117[15] = |(datain[251:248] ^ 3);
  assign w117[16] = |(datain[247:244] ^ 12);
  assign w117[17] = |(datain[243:240] ^ 0);
  assign w117[18] = |(datain[239:236] ^ 8);
  assign w117[19] = |(datain[235:232] ^ 14);
  assign w117[20] = |(datain[231:228] ^ 12);
  assign w117[21] = |(datain[227:224] ^ 0);
  assign w117[22] = |(datain[223:220] ^ 11);
  assign w117[23] = |(datain[219:216] ^ 8);
  assign w117[24] = |(datain[215:212] ^ 15);
  assign w117[25] = |(datain[211:208] ^ 0);
  assign w117[26] = |(datain[207:204] ^ 15);
  assign w117[27] = |(datain[203:200] ^ 0);
  assign w117[28] = |(datain[199:196] ^ 2);
  assign w117[29] = |(datain[195:192] ^ 6);
  assign comp[117] = ~(|w117);
  wire [32-1:0] w118;
  assign w118[0] = |(datain[311:308] ^ 0);
  assign w118[1] = |(datain[307:304] ^ 6);
  assign w118[2] = |(datain[303:300] ^ 0);
  assign w118[3] = |(datain[299:296] ^ 6);
  assign w118[4] = |(datain[295:292] ^ 0);
  assign w118[5] = |(datain[291:288] ^ 0);
  assign w118[6] = |(datain[287:284] ^ 5);
  assign w118[7] = |(datain[283:280] ^ 14);
  assign w118[8] = |(datain[279:276] ^ 5);
  assign w118[9] = |(datain[275:272] ^ 6);
  assign w118[10] = |(datain[271:268] ^ 1);
  assign w118[11] = |(datain[267:264] ^ 14);
  assign w118[12] = |(datain[263:260] ^ 0);
  assign w118[13] = |(datain[259:256] ^ 14);
  assign w118[14] = |(datain[255:252] ^ 3);
  assign w118[15] = |(datain[251:248] ^ 3);
  assign w118[16] = |(datain[247:244] ^ 15);
  assign w118[17] = |(datain[243:240] ^ 15);
  assign w118[18] = |(datain[239:236] ^ 8);
  assign w118[19] = |(datain[235:232] ^ 14);
  assign w118[20] = |(datain[231:228] ^ 13);
  assign w118[21] = |(datain[227:224] ^ 15);
  assign w118[22] = |(datain[223:220] ^ 12);
  assign w118[23] = |(datain[219:216] ^ 5);
  assign w118[24] = |(datain[215:212] ^ 0);
  assign w118[25] = |(datain[211:208] ^ 6);
  assign w118[26] = |(datain[207:204] ^ 8);
  assign w118[27] = |(datain[203:200] ^ 4);
  assign w118[28] = |(datain[199:196] ^ 0);
  assign w118[29] = |(datain[195:192] ^ 0);
  assign w118[30] = |(datain[191:188] ^ 2);
  assign w118[31] = |(datain[187:184] ^ 14);
  assign comp[118] = ~(|w118);
  wire [74-1:0] w119;
  assign w119[0] = |(datain[311:308] ^ 0);
  assign w119[1] = |(datain[307:304] ^ 5);
  assign w119[2] = |(datain[303:300] ^ 14);
  assign w119[3] = |(datain[299:296] ^ 9);
  assign w119[4] = |(datain[295:292] ^ 8);
  assign w119[5] = |(datain[291:288] ^ 0);
  assign w119[6] = |(datain[287:284] ^ 2);
  assign w119[7] = |(datain[283:280] ^ 14);
  assign w119[8] = |(datain[279:276] ^ 6);
  assign w119[9] = |(datain[275:272] ^ 10);
  assign w119[10] = |(datain[271:268] ^ 0);
  assign w119[11] = |(datain[267:264] ^ 5);
  assign w119[12] = |(datain[263:260] ^ 0);
  assign w119[13] = |(datain[259:256] ^ 3);
  assign w119[14] = |(datain[255:252] ^ 11);
  assign w119[15] = |(datain[251:248] ^ 4);
  assign w119[16] = |(datain[247:244] ^ 4);
  assign w119[17] = |(datain[243:240] ^ 0);
  assign w119[18] = |(datain[239:236] ^ 11);
  assign w119[19] = |(datain[235:232] ^ 9);
  assign w119[20] = |(datain[231:228] ^ 0);
  assign w119[21] = |(datain[227:224] ^ 3);
  assign w119[22] = |(datain[223:220] ^ 0);
  assign w119[23] = |(datain[219:216] ^ 0);
  assign w119[24] = |(datain[215:212] ^ 11);
  assign w119[25] = |(datain[211:208] ^ 10);
  assign w119[26] = |(datain[207:204] ^ 6);
  assign w119[27] = |(datain[203:200] ^ 9);
  assign w119[28] = |(datain[199:196] ^ 0);
  assign w119[29] = |(datain[195:192] ^ 5);
  assign w119[30] = |(datain[191:188] ^ 12);
  assign w119[31] = |(datain[187:184] ^ 13);
  assign w119[32] = |(datain[183:180] ^ 2);
  assign w119[33] = |(datain[179:176] ^ 1);
  assign w119[34] = |(datain[175:172] ^ 11);
  assign w119[35] = |(datain[171:168] ^ 0);
  assign w119[36] = |(datain[167:164] ^ 0);
  assign w119[37] = |(datain[163:160] ^ 2);
  assign w119[38] = |(datain[159:156] ^ 14);
  assign w119[39] = |(datain[155:152] ^ 8);
  assign w119[40] = |(datain[151:148] ^ 9);
  assign w119[41] = |(datain[147:144] ^ 13);
  assign w119[42] = |(datain[143:140] ^ 15);
  assign w119[43] = |(datain[139:136] ^ 15);
  assign w119[44] = |(datain[135:132] ^ 2);
  assign w119[45] = |(datain[131:128] ^ 13);
  assign w119[46] = |(datain[127:124] ^ 0);
  assign w119[47] = |(datain[123:120] ^ 7);
  assign w119[48] = |(datain[119:116] ^ 0);
  assign w119[49] = |(datain[115:112] ^ 0);
  assign w119[50] = |(datain[111:108] ^ 8);
  assign w119[51] = |(datain[107:104] ^ 11);
  assign w119[52] = |(datain[103:100] ^ 12);
  assign w119[53] = |(datain[99:96] ^ 10);
  assign w119[54] = |(datain[95:92] ^ 8);
  assign w119[55] = |(datain[91:88] ^ 11);
  assign w119[56] = |(datain[87:84] ^ 13);
  assign w119[57] = |(datain[83:80] ^ 0);
  assign w119[58] = |(datain[79:76] ^ 11);
  assign w119[59] = |(datain[75:72] ^ 8);
  assign w119[60] = |(datain[71:68] ^ 0);
  assign w119[61] = |(datain[67:64] ^ 0);
  assign w119[62] = |(datain[63:60] ^ 4);
  assign w119[63] = |(datain[59:56] ^ 2);
  assign w119[64] = |(datain[55:52] ^ 12);
  assign w119[65] = |(datain[51:48] ^ 13);
  assign w119[66] = |(datain[47:44] ^ 2);
  assign w119[67] = |(datain[43:40] ^ 1);
  assign w119[68] = |(datain[39:36] ^ 11);
  assign w119[69] = |(datain[35:32] ^ 4);
  assign w119[70] = |(datain[31:28] ^ 3);
  assign w119[71] = |(datain[27:24] ^ 15);
  assign w119[72] = |(datain[23:20] ^ 11);
  assign w119[73] = |(datain[19:16] ^ 9);
  assign comp[119] = ~(|w119);
  wire [76-1:0] w120;
  assign w120[0] = |(datain[311:308] ^ 0);
  assign w120[1] = |(datain[307:304] ^ 2);
  assign w120[2] = |(datain[303:300] ^ 3);
  assign w120[3] = |(datain[299:296] ^ 13);
  assign w120[4] = |(datain[295:292] ^ 11);
  assign w120[5] = |(datain[291:288] ^ 10);
  assign w120[6] = |(datain[287:284] ^ 9);
  assign w120[7] = |(datain[283:280] ^ 14);
  assign w120[8] = |(datain[279:276] ^ 0);
  assign w120[9] = |(datain[275:272] ^ 0);
  assign w120[10] = |(datain[271:268] ^ 12);
  assign w120[11] = |(datain[267:264] ^ 13);
  assign w120[12] = |(datain[263:260] ^ 2);
  assign w120[13] = |(datain[259:256] ^ 1);
  assign w120[14] = |(datain[255:252] ^ 9);
  assign w120[15] = |(datain[251:248] ^ 3);
  assign w120[16] = |(datain[247:244] ^ 11);
  assign w120[17] = |(datain[243:240] ^ 9);
  assign w120[18] = |(datain[239:236] ^ 1);
  assign w120[19] = |(datain[235:232] ^ 1);
  assign w120[20] = |(datain[231:228] ^ 0);
  assign w120[21] = |(datain[227:224] ^ 3);
  assign w120[22] = |(datain[223:220] ^ 11);
  assign w120[23] = |(datain[219:216] ^ 4);
  assign w120[24] = |(datain[215:212] ^ 4);
  assign w120[25] = |(datain[211:208] ^ 0);
  assign w120[26] = |(datain[207:204] ^ 11);
  assign w120[27] = |(datain[203:200] ^ 10);
  assign w120[28] = |(datain[199:196] ^ 0);
  assign w120[29] = |(datain[195:192] ^ 0);
  assign w120[30] = |(datain[191:188] ^ 0);
  assign w120[31] = |(datain[187:184] ^ 1);
  assign w120[32] = |(datain[183:180] ^ 12);
  assign w120[33] = |(datain[179:176] ^ 13);
  assign w120[34] = |(datain[175:172] ^ 2);
  assign w120[35] = |(datain[171:168] ^ 1);
  assign w120[36] = |(datain[167:164] ^ 11);
  assign w120[37] = |(datain[163:160] ^ 4);
  assign w120[38] = |(datain[159:156] ^ 3);
  assign w120[39] = |(datain[155:152] ^ 14);
  assign w120[40] = |(datain[151:148] ^ 12);
  assign w120[41] = |(datain[147:144] ^ 13);
  assign w120[42] = |(datain[143:140] ^ 2);
  assign w120[43] = |(datain[139:136] ^ 1);
  assign w120[44] = |(datain[135:132] ^ 15);
  assign w120[45] = |(datain[131:128] ^ 15);
  assign w120[46] = |(datain[127:124] ^ 0);
  assign w120[47] = |(datain[123:120] ^ 6);
  assign w120[48] = |(datain[119:116] ^ 0);
  assign w120[49] = |(datain[115:112] ^ 12);
  assign w120[50] = |(datain[111:108] ^ 0);
  assign w120[51] = |(datain[107:104] ^ 4);
  assign w120[52] = |(datain[103:100] ^ 8);
  assign w120[53] = |(datain[99:96] ^ 3);
  assign w120[54] = |(datain[95:92] ^ 3);
  assign w120[55] = |(datain[91:88] ^ 14);
  assign w120[56] = |(datain[87:84] ^ 0);
  assign w120[57] = |(datain[83:80] ^ 12);
  assign w120[58] = |(datain[79:76] ^ 0);
  assign w120[59] = |(datain[75:72] ^ 4);
  assign w120[60] = |(datain[71:68] ^ 0);
  assign w120[61] = |(datain[67:64] ^ 5);
  assign w120[62] = |(datain[63:60] ^ 7);
  assign w120[63] = |(datain[59:56] ^ 13);
  assign w120[64] = |(datain[55:52] ^ 0);
  assign w120[65] = |(datain[51:48] ^ 3);
  assign w120[66] = |(datain[47:44] ^ 14);
  assign w120[67] = |(datain[43:40] ^ 8);
  assign w120[68] = |(datain[39:36] ^ 13);
  assign w120[69] = |(datain[35:32] ^ 4);
  assign w120[70] = |(datain[31:28] ^ 15);
  assign w120[71] = |(datain[27:24] ^ 15);
  assign w120[72] = |(datain[23:20] ^ 11);
  assign w120[73] = |(datain[19:16] ^ 4);
  assign w120[74] = |(datain[15:12] ^ 3);
  assign w120[75] = |(datain[11:8] ^ 11);
  assign comp[120] = ~(|w120);
  wire [32-1:0] w121;
  assign w121[0] = |(datain[311:308] ^ 0);
  assign w121[1] = |(datain[307:304] ^ 1);
  assign w121[2] = |(datain[303:300] ^ 8);
  assign w121[3] = |(datain[299:296] ^ 10);
  assign w121[4] = |(datain[295:292] ^ 5);
  assign w121[5] = |(datain[291:288] ^ 4);
  assign w121[6] = |(datain[287:284] ^ 0);
  assign w121[7] = |(datain[283:280] ^ 5);
  assign w121[8] = |(datain[279:276] ^ 8);
  assign w121[9] = |(datain[275:272] ^ 8);
  assign w121[10] = |(datain[271:268] ^ 1);
  assign w121[11] = |(datain[267:264] ^ 6);
  assign w121[12] = |(datain[263:260] ^ 0);
  assign w121[13] = |(datain[259:256] ^ 0);
  assign w121[14] = |(datain[255:252] ^ 0);
  assign w121[15] = |(datain[251:248] ^ 1);
  assign w121[16] = |(datain[247:244] ^ 11);
  assign w121[17] = |(datain[243:240] ^ 4);
  assign w121[18] = |(datain[239:236] ^ 2);
  assign w121[19] = |(datain[235:232] ^ 10);
  assign w121[20] = |(datain[231:228] ^ 12);
  assign w121[21] = |(datain[227:224] ^ 13);
  assign w121[22] = |(datain[223:220] ^ 2);
  assign w121[23] = |(datain[219:216] ^ 1);
  assign w121[24] = |(datain[215:212] ^ 15);
  assign w121[25] = |(datain[211:208] ^ 6);
  assign w121[26] = |(datain[207:204] ^ 12);
  assign w121[27] = |(datain[203:200] ^ 2);
  assign w121[28] = |(datain[199:196] ^ 0);
  assign w121[29] = |(datain[195:192] ^ 1);
  assign w121[30] = |(datain[191:188] ^ 7);
  assign w121[31] = |(datain[187:184] ^ 5);
  assign comp[121] = ~(|w121);
  wire [36-1:0] w122;
  assign w122[0] = |(datain[311:308] ^ 0);
  assign w122[1] = |(datain[307:304] ^ 2);
  assign w122[2] = |(datain[303:300] ^ 4);
  assign w122[3] = |(datain[299:296] ^ 2);
  assign w122[4] = |(datain[295:292] ^ 14);
  assign w122[5] = |(datain[291:288] ^ 8);
  assign w122[6] = |(datain[287:284] ^ 8);
  assign w122[7] = |(datain[283:280] ^ 12);
  assign w122[8] = |(datain[279:276] ^ 0);
  assign w122[9] = |(datain[275:272] ^ 0);
  assign w122[10] = |(datain[271:268] ^ 11);
  assign w122[11] = |(datain[267:264] ^ 4);
  assign w122[12] = |(datain[263:260] ^ 4);
  assign w122[13] = |(datain[259:256] ^ 0);
  assign w122[14] = |(datain[255:252] ^ 11);
  assign w122[15] = |(datain[251:248] ^ 9);
  assign w122[16] = |(datain[247:244] ^ 2);
  assign w122[17] = |(datain[243:240] ^ 11);
  assign w122[18] = |(datain[239:236] ^ 0);
  assign w122[19] = |(datain[235:232] ^ 4);
  assign w122[20] = |(datain[231:228] ^ 9);
  assign w122[21] = |(datain[227:224] ^ 0);
  assign w122[22] = |(datain[223:220] ^ 11);
  assign w122[23] = |(datain[219:216] ^ 10);
  assign w122[24] = |(datain[215:212] ^ 0);
  assign w122[25] = |(datain[211:208] ^ 0);
  assign w122[26] = |(datain[207:204] ^ 0);
  assign w122[27] = |(datain[203:200] ^ 1);
  assign w122[28] = |(datain[199:196] ^ 12);
  assign w122[29] = |(datain[195:192] ^ 13);
  assign w122[30] = |(datain[191:188] ^ 2);
  assign w122[31] = |(datain[187:184] ^ 1);
  assign w122[32] = |(datain[183:180] ^ 7);
  assign w122[33] = |(datain[179:176] ^ 2);
  assign w122[34] = |(datain[175:172] ^ 1);
  assign w122[35] = |(datain[171:168] ^ 4);
  assign comp[122] = ~(|w122);
  wire [32-1:0] w123;
  assign w123[0] = |(datain[311:308] ^ 4);
  assign w123[1] = |(datain[307:304] ^ 14);
  assign w123[2] = |(datain[303:300] ^ 0);
  assign w123[3] = |(datain[299:296] ^ 1);
  assign w123[4] = |(datain[295:292] ^ 14);
  assign w123[5] = |(datain[291:288] ^ 10);
  assign w123[6] = |(datain[287:284] ^ 12);
  assign w123[7] = |(datain[283:280] ^ 13);
  assign w123[8] = |(datain[279:276] ^ 2);
  assign w123[9] = |(datain[275:272] ^ 1);
  assign w123[10] = |(datain[271:268] ^ 12);
  assign w123[11] = |(datain[267:264] ^ 3);
  assign w123[12] = |(datain[263:260] ^ 11);
  assign w123[13] = |(datain[259:256] ^ 4);
  assign w123[14] = |(datain[255:252] ^ 4);
  assign w123[15] = |(datain[251:248] ^ 15);
  assign w123[16] = |(datain[247:244] ^ 12);
  assign w123[17] = |(datain[243:240] ^ 13);
  assign w123[18] = |(datain[239:236] ^ 2);
  assign w123[19] = |(datain[235:232] ^ 1);
  assign w123[20] = |(datain[231:228] ^ 12);
  assign w123[21] = |(datain[227:224] ^ 3);
  assign w123[22] = |(datain[223:220] ^ 5);
  assign w123[23] = |(datain[219:216] ^ 1);
  assign w123[24] = |(datain[215:212] ^ 3);
  assign w123[25] = |(datain[211:208] ^ 3);
  assign w123[26] = |(datain[207:204] ^ 12);
  assign w123[27] = |(datain[203:200] ^ 0);
  assign w123[28] = |(datain[199:196] ^ 3);
  assign w123[29] = |(datain[195:192] ^ 11);
  assign w123[30] = |(datain[191:188] ^ 8);
  assign w123[31] = |(datain[187:184] ^ 6);
  assign comp[123] = ~(|w123);
  wire [30-1:0] w124;
  assign w124[0] = |(datain[311:308] ^ 4);
  assign w124[1] = |(datain[307:304] ^ 0);
  assign w124[2] = |(datain[303:300] ^ 0);
  assign w124[3] = |(datain[299:296] ^ 0);
  assign w124[4] = |(datain[295:292] ^ 8);
  assign w124[5] = |(datain[291:288] ^ 14);
  assign w124[6] = |(datain[287:284] ^ 13);
  assign w124[7] = |(datain[283:280] ^ 8);
  assign w124[8] = |(datain[279:276] ^ 10);
  assign w124[9] = |(datain[275:272] ^ 1);
  assign w124[10] = |(datain[271:268] ^ 1);
  assign w124[11] = |(datain[267:264] ^ 3);
  assign w124[12] = |(datain[263:260] ^ 0);
  assign w124[13] = |(datain[259:256] ^ 0);
  assign w124[14] = |(datain[255:252] ^ 11);
  assign w124[15] = |(datain[251:248] ^ 1);
  assign w124[16] = |(datain[247:244] ^ 0);
  assign w124[17] = |(datain[243:240] ^ 6);
  assign w124[18] = |(datain[239:236] ^ 13);
  assign w124[19] = |(datain[235:232] ^ 3);
  assign w124[20] = |(datain[231:228] ^ 14);
  assign w124[21] = |(datain[227:224] ^ 0);
  assign w124[22] = |(datain[223:220] ^ 2);
  assign w124[23] = |(datain[219:216] ^ 13);
  assign w124[24] = |(datain[215:212] ^ 0);
  assign w124[25] = |(datain[211:208] ^ 0);
  assign w124[26] = |(datain[207:204] ^ 0);
  assign w124[27] = |(datain[203:200] ^ 8);
  assign w124[28] = |(datain[199:196] ^ 8);
  assign w124[29] = |(datain[195:192] ^ 14);
  assign comp[124] = ~(|w124);
  wire [38-1:0] w125;
  assign w125[0] = |(datain[311:308] ^ 0);
  assign w125[1] = |(datain[307:304] ^ 1);
  assign w125[2] = |(datain[303:300] ^ 7);
  assign w125[3] = |(datain[299:296] ^ 5);
  assign w125[4] = |(datain[295:292] ^ 13);
  assign w125[5] = |(datain[291:288] ^ 0);
  assign w125[6] = |(datain[287:284] ^ 0);
  assign w125[7] = |(datain[283:280] ^ 14);
  assign w125[8] = |(datain[279:276] ^ 0);
  assign w125[9] = |(datain[275:272] ^ 14);
  assign w125[10] = |(datain[271:268] ^ 1);
  assign w125[11] = |(datain[267:264] ^ 15);
  assign w125[12] = |(datain[263:260] ^ 0);
  assign w125[13] = |(datain[259:256] ^ 7);
  assign w125[14] = |(datain[255:252] ^ 11);
  assign w125[15] = |(datain[251:248] ^ 14);
  assign w125[16] = |(datain[247:244] ^ 13);
  assign w125[17] = |(datain[243:240] ^ 3);
  assign w125[18] = |(datain[239:236] ^ 0);
  assign w125[19] = |(datain[235:232] ^ 4);
  assign w125[20] = |(datain[231:228] ^ 2);
  assign w125[21] = |(datain[227:224] ^ 11);
  assign w125[22] = |(datain[223:220] ^ 12);
  assign w125[23] = |(datain[219:216] ^ 9);
  assign w125[24] = |(datain[215:212] ^ 2);
  assign w125[25] = |(datain[211:208] ^ 14);
  assign w125[26] = |(datain[207:204] ^ 8);
  assign w125[27] = |(datain[203:200] ^ 10);
  assign w125[28] = |(datain[199:196] ^ 0);
  assign w125[29] = |(datain[195:192] ^ 4);
  assign w125[30] = |(datain[191:188] ^ 4);
  assign w125[31] = |(datain[187:184] ^ 6);
  assign w125[32] = |(datain[183:180] ^ 4);
  assign w125[33] = |(datain[179:176] ^ 1);
  assign w125[34] = |(datain[175:172] ^ 0);
  assign w125[35] = |(datain[171:168] ^ 10);
  assign w125[36] = |(datain[167:164] ^ 12);
  assign w125[37] = |(datain[163:160] ^ 0);
  assign comp[125] = ~(|w125);
  wire [30-1:0] w126;
  assign w126[0] = |(datain[311:308] ^ 11);
  assign w126[1] = |(datain[307:304] ^ 15);
  assign w126[2] = |(datain[303:300] ^ 0);
  assign w126[3] = |(datain[299:296] ^ 0);
  assign w126[4] = |(datain[295:292] ^ 0);
  assign w126[5] = |(datain[291:288] ^ 1);
  assign w126[6] = |(datain[287:284] ^ 4);
  assign w126[7] = |(datain[283:280] ^ 7);
  assign w126[8] = |(datain[279:276] ^ 0);
  assign w126[9] = |(datain[275:272] ^ 3);
  assign w126[10] = |(datain[271:268] ^ 3);
  assign w126[11] = |(datain[267:264] ^ 13);
  assign w126[12] = |(datain[263:260] ^ 8);
  assign w126[13] = |(datain[259:256] ^ 11);
  assign w126[14] = |(datain[255:252] ^ 15);
  assign w126[15] = |(datain[251:248] ^ 7);
  assign w126[16] = |(datain[247:244] ^ 3);
  assign w126[17] = |(datain[243:240] ^ 3);
  assign w126[18] = |(datain[239:236] ^ 12);
  assign w126[19] = |(datain[235:232] ^ 0);
  assign w126[20] = |(datain[231:228] ^ 11);
  assign w126[21] = |(datain[227:224] ^ 10);
  assign w126[22] = |(datain[223:220] ^ 5);
  assign w126[23] = |(datain[219:216] ^ 4);
  assign w126[24] = |(datain[215:212] ^ 0);
  assign w126[25] = |(datain[211:208] ^ 2);
  assign w126[26] = |(datain[207:204] ^ 5);
  assign w126[27] = |(datain[203:200] ^ 2);
  assign w126[28] = |(datain[199:196] ^ 3);
  assign w126[29] = |(datain[195:192] ^ 3);
  assign comp[126] = ~(|w126);
  wire [44-1:0] w127;
  assign w127[0] = |(datain[311:308] ^ 0);
  assign w127[1] = |(datain[307:304] ^ 3);
  assign w127[2] = |(datain[303:300] ^ 11);
  assign w127[3] = |(datain[299:296] ^ 15);
  assign w127[4] = |(datain[295:292] ^ 0);
  assign w127[5] = |(datain[291:288] ^ 0);
  assign w127[6] = |(datain[287:284] ^ 0);
  assign w127[7] = |(datain[283:280] ^ 9);
  assign w127[8] = |(datain[279:276] ^ 14);
  assign w127[9] = |(datain[275:272] ^ 8);
  assign w127[10] = |(datain[271:268] ^ 1);
  assign w127[11] = |(datain[267:264] ^ 14);
  assign w127[12] = |(datain[263:260] ^ 15);
  assign w127[13] = |(datain[259:256] ^ 15);
  assign w127[14] = |(datain[255:252] ^ 14);
  assign w127[15] = |(datain[251:248] ^ 8);
  assign w127[16] = |(datain[247:244] ^ 1);
  assign w127[17] = |(datain[243:240] ^ 11);
  assign w127[18] = |(datain[239:236] ^ 15);
  assign w127[19] = |(datain[235:232] ^ 15);
  assign w127[20] = |(datain[231:228] ^ 11);
  assign w127[21] = |(datain[227:224] ^ 11);
  assign w127[22] = |(datain[223:220] ^ 3);
  assign w127[23] = |(datain[219:216] ^ 15);
  assign w127[24] = |(datain[215:212] ^ 0);
  assign w127[25] = |(datain[211:208] ^ 0);
  assign w127[26] = |(datain[207:204] ^ 11);
  assign w127[27] = |(datain[203:200] ^ 10);
  assign w127[28] = |(datain[199:196] ^ 15);
  assign w127[29] = |(datain[195:192] ^ 15);
  assign w127[30] = |(datain[191:188] ^ 0);
  assign w127[31] = |(datain[187:184] ^ 0);
  assign w127[32] = |(datain[183:180] ^ 8);
  assign w127[33] = |(datain[179:176] ^ 10);
  assign w127[34] = |(datain[175:172] ^ 12);
  assign w127[35] = |(datain[171:168] ^ 3);
  assign w127[36] = |(datain[167:164] ^ 8);
  assign w127[37] = |(datain[163:160] ^ 11);
  assign w127[38] = |(datain[159:156] ^ 15);
  assign w127[39] = |(datain[155:152] ^ 3);
  assign w127[40] = |(datain[151:148] ^ 8);
  assign w127[41] = |(datain[147:144] ^ 11);
  assign w127[42] = |(datain[143:140] ^ 11);
  assign w127[43] = |(datain[139:136] ^ 0);
  assign comp[127] = ~(|w127);
  wire [32-1:0] w128;
  assign w128[0] = |(datain[311:308] ^ 8);
  assign w128[1] = |(datain[307:304] ^ 10);
  assign w128[2] = |(datain[303:300] ^ 4);
  assign w128[3] = |(datain[299:296] ^ 6);
  assign w128[4] = |(datain[295:292] ^ 0);
  assign w128[5] = |(datain[291:288] ^ 0);
  assign w128[6] = |(datain[287:284] ^ 10);
  assign w128[7] = |(datain[283:280] ^ 2);
  assign w128[8] = |(datain[279:276] ^ 0);
  assign w128[9] = |(datain[275:272] ^ 0);
  assign w128[10] = |(datain[271:268] ^ 0);
  assign w128[11] = |(datain[267:264] ^ 1);
  assign w128[12] = |(datain[263:260] ^ 8);
  assign w128[13] = |(datain[259:256] ^ 11);
  assign w128[14] = |(datain[255:252] ^ 4);
  assign w128[15] = |(datain[251:248] ^ 6);
  assign w128[16] = |(datain[247:244] ^ 0);
  assign w128[17] = |(datain[243:240] ^ 1);
  assign w128[18] = |(datain[239:236] ^ 10);
  assign w128[19] = |(datain[235:232] ^ 3);
  assign w128[20] = |(datain[231:228] ^ 0);
  assign w128[21] = |(datain[227:224] ^ 1);
  assign w128[22] = |(datain[223:220] ^ 0);
  assign w128[23] = |(datain[219:216] ^ 1);
  assign w128[24] = |(datain[215:212] ^ 11);
  assign w128[25] = |(datain[211:208] ^ 8);
  assign w128[26] = |(datain[207:204] ^ 12);
  assign w128[27] = |(datain[203:200] ^ 12);
  assign w128[28] = |(datain[199:196] ^ 4);
  assign w128[29] = |(datain[195:192] ^ 11);
  assign w128[30] = |(datain[191:188] ^ 12);
  assign w128[31] = |(datain[187:184] ^ 13);
  assign comp[128] = ~(|w128);
  wire [32-1:0] w129;
  assign w129[0] = |(datain[311:308] ^ 12);
  assign w129[1] = |(datain[307:304] ^ 13);
  assign w129[2] = |(datain[303:300] ^ 2);
  assign w129[3] = |(datain[299:296] ^ 1);
  assign w129[4] = |(datain[295:292] ^ 7);
  assign w129[5] = |(datain[291:288] ^ 2);
  assign w129[6] = |(datain[287:284] ^ 5);
  assign w129[7] = |(datain[283:280] ^ 2);
  assign w129[8] = |(datain[279:276] ^ 11);
  assign w129[9] = |(datain[275:272] ^ 9);
  assign w129[10] = |(datain[271:268] ^ 1);
  assign w129[11] = |(datain[267:264] ^ 14);
  assign w129[12] = |(datain[263:260] ^ 0);
  assign w129[13] = |(datain[259:256] ^ 0);
  assign w129[14] = |(datain[255:252] ^ 11);
  assign w129[15] = |(datain[251:248] ^ 10);
  assign w129[16] = |(datain[247:244] ^ 7);
  assign w129[17] = |(datain[243:240] ^ 13);
  assign w129[18] = |(datain[239:236] ^ 0);
  assign w129[19] = |(datain[235:232] ^ 4);
  assign w129[20] = |(datain[231:228] ^ 11);
  assign w129[21] = |(datain[227:224] ^ 4);
  assign w129[22] = |(datain[223:220] ^ 3);
  assign w129[23] = |(datain[219:216] ^ 15);
  assign w129[24] = |(datain[215:212] ^ 12);
  assign w129[25] = |(datain[211:208] ^ 13);
  assign w129[26] = |(datain[207:204] ^ 2);
  assign w129[27] = |(datain[203:200] ^ 1);
  assign w129[28] = |(datain[199:196] ^ 7);
  assign w129[29] = |(datain[195:192] ^ 2);
  assign w129[30] = |(datain[191:188] ^ 4);
  assign w129[31] = |(datain[187:184] ^ 6);
  assign comp[129] = ~(|w129);
  wire [76-1:0] w130;
  assign w130[0] = |(datain[311:308] ^ 11);
  assign w130[1] = |(datain[307:304] ^ 9);
  assign w130[2] = |(datain[303:300] ^ 3);
  assign w130[3] = |(datain[299:296] ^ 14);
  assign w130[4] = |(datain[295:292] ^ 0);
  assign w130[5] = |(datain[291:288] ^ 0);
  assign w130[6] = |(datain[287:284] ^ 11);
  assign w130[7] = |(datain[283:280] ^ 10);
  assign w130[8] = |(datain[279:276] ^ 12);
  assign w130[9] = |(datain[275:272] ^ 9);
  assign w130[10] = |(datain[271:268] ^ 0);
  assign w130[11] = |(datain[267:264] ^ 9);
  assign w130[12] = |(datain[263:260] ^ 14);
  assign w130[13] = |(datain[259:256] ^ 11);
  assign w130[14] = |(datain[255:252] ^ 0);
  assign w130[15] = |(datain[251:248] ^ 6);
  assign w130[16] = |(datain[247:244] ^ 11);
  assign w130[17] = |(datain[243:240] ^ 9);
  assign w130[18] = |(datain[239:236] ^ 1);
  assign w130[19] = |(datain[235:232] ^ 13);
  assign w130[20] = |(datain[231:228] ^ 0);
  assign w130[21] = |(datain[227:224] ^ 0);
  assign w130[22] = |(datain[223:220] ^ 11);
  assign w130[23] = |(datain[219:216] ^ 10);
  assign w130[24] = |(datain[215:212] ^ 0);
  assign w130[25] = |(datain[211:208] ^ 7);
  assign w130[26] = |(datain[207:204] ^ 0);
  assign w130[27] = |(datain[203:200] ^ 10);
  assign w130[28] = |(datain[199:196] ^ 11);
  assign w130[29] = |(datain[195:192] ^ 4);
  assign w130[30] = |(datain[191:188] ^ 4);
  assign w130[31] = |(datain[187:184] ^ 0);
  assign w130[32] = |(datain[183:180] ^ 12);
  assign w130[33] = |(datain[179:176] ^ 13);
  assign w130[34] = |(datain[175:172] ^ 2);
  assign w130[35] = |(datain[171:168] ^ 1);
  assign w130[36] = |(datain[167:164] ^ 11);
  assign w130[37] = |(datain[163:160] ^ 8);
  assign w130[38] = |(datain[159:156] ^ 0);
  assign w130[39] = |(datain[155:152] ^ 0);
  assign w130[40] = |(datain[151:148] ^ 4);
  assign w130[41] = |(datain[147:144] ^ 2);
  assign w130[42] = |(datain[143:140] ^ 3);
  assign w130[43] = |(datain[139:136] ^ 3);
  assign w130[44] = |(datain[135:132] ^ 12);
  assign w130[45] = |(datain[131:128] ^ 9);
  assign w130[46] = |(datain[127:124] ^ 9);
  assign w130[47] = |(datain[123:120] ^ 9);
  assign w130[48] = |(datain[119:116] ^ 12);
  assign w130[49] = |(datain[115:112] ^ 13);
  assign w130[50] = |(datain[111:108] ^ 2);
  assign w130[51] = |(datain[107:104] ^ 1);
  assign w130[52] = |(datain[103:100] ^ 11);
  assign w130[53] = |(datain[99:96] ^ 4);
  assign w130[54] = |(datain[95:92] ^ 4);
  assign w130[55] = |(datain[91:88] ^ 0);
  assign w130[56] = |(datain[87:84] ^ 11);
  assign w130[57] = |(datain[83:80] ^ 9);
  assign w130[58] = |(datain[79:76] ^ 5);
  assign w130[59] = |(datain[75:72] ^ 10);
  assign w130[60] = |(datain[71:68] ^ 0);
  assign w130[61] = |(datain[67:64] ^ 0);
  assign w130[62] = |(datain[63:60] ^ 11);
  assign w130[63] = |(datain[59:56] ^ 10);
  assign w130[64] = |(datain[55:52] ^ 4);
  assign w130[65] = |(datain[51:48] ^ 6);
  assign w130[66] = |(datain[47:44] ^ 0);
  assign w130[67] = |(datain[43:40] ^ 8);
  assign w130[68] = |(datain[39:36] ^ 12);
  assign w130[69] = |(datain[35:32] ^ 13);
  assign w130[70] = |(datain[31:28] ^ 2);
  assign w130[71] = |(datain[27:24] ^ 1);
  assign w130[72] = |(datain[23:20] ^ 12);
  assign w130[73] = |(datain[19:16] ^ 3);
  assign w130[74] = |(datain[15:12] ^ 10);
  assign w130[75] = |(datain[11:8] ^ 1);
  assign comp[130] = ~(|w130);
  wire [28-1:0] w131;
  assign w131[0] = |(datain[311:308] ^ 8);
  assign w131[1] = |(datain[307:304] ^ 12);
  assign w131[2] = |(datain[303:300] ^ 12);
  assign w131[3] = |(datain[299:296] ^ 8);
  assign w131[4] = |(datain[295:292] ^ 8);
  assign w131[5] = |(datain[291:288] ^ 14);
  assign w131[6] = |(datain[287:284] ^ 13);
  assign w131[7] = |(datain[283:280] ^ 0);
  assign w131[8] = |(datain[279:276] ^ 11);
  assign w131[9] = |(datain[275:272] ^ 12);
  assign w131[10] = |(datain[271:268] ^ 0);
  assign w131[11] = |(datain[267:264] ^ 0);
  assign w131[12] = |(datain[263:260] ^ 7);
  assign w131[13] = |(datain[259:256] ^ 12);
  assign w131[14] = |(datain[255:252] ^ 8);
  assign w131[15] = |(datain[251:248] ^ 11);
  assign w131[16] = |(datain[247:244] ^ 15);
  assign w131[17] = |(datain[243:240] ^ 4);
  assign w131[18] = |(datain[239:236] ^ 8);
  assign w131[19] = |(datain[235:232] ^ 14);
  assign w131[20] = |(datain[231:228] ^ 12);
  assign w131[21] = |(datain[227:224] ^ 0);
  assign w131[22] = |(datain[223:220] ^ 8);
  assign w131[23] = |(datain[219:216] ^ 14);
  assign w131[24] = |(datain[215:212] ^ 13);
  assign w131[25] = |(datain[211:208] ^ 8);
  assign w131[26] = |(datain[207:204] ^ 5);
  assign w131[27] = |(datain[203:200] ^ 0);
  assign comp[131] = ~(|w131);
  wire [74-1:0] w132;
  assign w132[0] = |(datain[311:308] ^ 4);
  assign w132[1] = |(datain[307:304] ^ 5);
  assign w132[2] = |(datain[303:300] ^ 1);
  assign w132[3] = |(datain[299:296] ^ 5);
  assign w132[4] = |(datain[295:292] ^ 0);
  assign w132[5] = |(datain[291:288] ^ 0);
  assign w132[6] = |(datain[287:284] ^ 0);
  assign w132[7] = |(datain[283:280] ^ 0);
  assign w132[8] = |(datain[279:276] ^ 2);
  assign w132[9] = |(datain[275:272] ^ 6);
  assign w132[10] = |(datain[271:268] ^ 12);
  assign w132[11] = |(datain[267:264] ^ 7);
  assign w132[12] = |(datain[263:260] ^ 4);
  assign w132[13] = |(datain[259:256] ^ 5);
  assign w132[14] = |(datain[255:252] ^ 1);
  assign w132[15] = |(datain[251:248] ^ 7);
  assign w132[16] = |(datain[247:244] ^ 0);
  assign w132[17] = |(datain[243:240] ^ 0);
  assign w132[18] = |(datain[239:236] ^ 0);
  assign w132[19] = |(datain[235:232] ^ 0);
  assign w132[20] = |(datain[231:228] ^ 11);
  assign w132[21] = |(datain[227:224] ^ 10);
  assign w132[22] = |(datain[223:220] ^ 15);
  assign w132[23] = |(datain[219:216] ^ 11);
  assign w132[24] = |(datain[215:212] ^ 0);
  assign w132[25] = |(datain[211:208] ^ 6);
  assign w132[26] = |(datain[207:204] ^ 11);
  assign w132[27] = |(datain[203:200] ^ 4);
  assign w132[28] = |(datain[199:196] ^ 4);
  assign w132[29] = |(datain[195:192] ^ 0);
  assign w132[30] = |(datain[191:188] ^ 12);
  assign w132[31] = |(datain[187:184] ^ 13);
  assign w132[32] = |(datain[183:180] ^ 2);
  assign w132[33] = |(datain[179:176] ^ 1);
  assign w132[34] = |(datain[175:172] ^ 2);
  assign w132[35] = |(datain[171:168] ^ 6);
  assign w132[36] = |(datain[167:164] ^ 8);
  assign w132[37] = |(datain[163:160] ^ 11);
  assign w132[38] = |(datain[159:156] ^ 4);
  assign w132[39] = |(datain[155:152] ^ 13);
  assign w132[40] = |(datain[151:148] ^ 0);
  assign w132[41] = |(datain[147:144] ^ 13);
  assign w132[42] = |(datain[143:140] ^ 2);
  assign w132[43] = |(datain[139:136] ^ 6);
  assign w132[44] = |(datain[135:132] ^ 8);
  assign w132[45] = |(datain[131:128] ^ 11);
  assign w132[46] = |(datain[127:124] ^ 5);
  assign w132[47] = |(datain[123:120] ^ 5);
  assign w132[48] = |(datain[119:116] ^ 0);
  assign w132[49] = |(datain[115:112] ^ 15);
  assign w132[50] = |(datain[111:108] ^ 13);
  assign w132[51] = |(datain[107:104] ^ 0);
  assign w132[52] = |(datain[103:100] ^ 12);
  assign w132[53] = |(datain[99:96] ^ 14);
  assign w132[54] = |(datain[95:92] ^ 8);
  assign w132[55] = |(datain[91:88] ^ 0);
  assign w132[56] = |(datain[87:84] ^ 12);
  assign w132[57] = |(datain[83:80] ^ 6);
  assign w132[58] = |(datain[79:76] ^ 6);
  assign w132[59] = |(datain[75:72] ^ 4);
  assign w132[60] = |(datain[71:68] ^ 13);
  assign w132[61] = |(datain[67:64] ^ 0);
  assign w132[62] = |(datain[63:60] ^ 12);
  assign w132[63] = |(datain[59:56] ^ 6);
  assign w132[64] = |(datain[55:52] ^ 11);
  assign w132[65] = |(datain[51:48] ^ 8);
  assign w132[66] = |(datain[47:44] ^ 0);
  assign w132[67] = |(datain[43:40] ^ 1);
  assign w132[68] = |(datain[39:36] ^ 5);
  assign w132[69] = |(datain[35:32] ^ 7);
  assign w132[70] = |(datain[31:28] ^ 12);
  assign w132[71] = |(datain[27:24] ^ 13);
  assign w132[72] = |(datain[23:20] ^ 2);
  assign w132[73] = |(datain[19:16] ^ 1);
  assign comp[132] = ~(|w132);
  wire [76-1:0] w133;
  assign w133[0] = |(datain[311:308] ^ 12);
  assign w133[1] = |(datain[307:304] ^ 3);
  assign w133[2] = |(datain[303:300] ^ 14);
  assign w133[3] = |(datain[299:296] ^ 8);
  assign w133[4] = |(datain[295:292] ^ 4);
  assign w133[5] = |(datain[291:288] ^ 6);
  assign w133[6] = |(datain[287:284] ^ 0);
  assign w133[7] = |(datain[283:280] ^ 0);
  assign w133[8] = |(datain[279:276] ^ 5);
  assign w133[9] = |(datain[275:272] ^ 11);
  assign w133[10] = |(datain[271:268] ^ 5);
  assign w133[11] = |(datain[267:264] ^ 15);
  assign w133[12] = |(datain[263:260] ^ 0);
  assign w133[13] = |(datain[259:256] ^ 7);
  assign w133[14] = |(datain[255:252] ^ 11);
  assign w133[15] = |(datain[251:248] ^ 4);
  assign w133[16] = |(datain[247:244] ^ 4);
  assign w133[17] = |(datain[243:240] ^ 0);
  assign w133[18] = |(datain[239:236] ^ 11);
  assign w133[19] = |(datain[235:232] ^ 9);
  assign w133[20] = |(datain[231:228] ^ 13);
  assign w133[21] = |(datain[227:224] ^ 10);
  assign w133[22] = |(datain[223:220] ^ 0);
  assign w133[23] = |(datain[219:216] ^ 5);
  assign w133[24] = |(datain[215:212] ^ 9);
  assign w133[25] = |(datain[211:208] ^ 0);
  assign w133[26] = |(datain[207:204] ^ 11);
  assign w133[27] = |(datain[203:200] ^ 10);
  assign w133[28] = |(datain[199:196] ^ 3);
  assign w133[29] = |(datain[195:192] ^ 3);
  assign w133[30] = |(datain[191:188] ^ 0);
  assign w133[31] = |(datain[187:184] ^ 7);
  assign w133[32] = |(datain[183:180] ^ 12);
  assign w133[33] = |(datain[179:176] ^ 13);
  assign w133[34] = |(datain[175:172] ^ 2);
  assign w133[35] = |(datain[171:168] ^ 1);
  assign w133[36] = |(datain[167:164] ^ 12);
  assign w133[37] = |(datain[163:160] ^ 3);
  assign w133[38] = |(datain[159:156] ^ 2);
  assign w133[39] = |(datain[155:152] ^ 6);
  assign w133[40] = |(datain[151:148] ^ 8);
  assign w133[41] = |(datain[147:144] ^ 11);
  assign w133[42] = |(datain[143:140] ^ 4);
  assign w133[43] = |(datain[139:136] ^ 5);
  assign w133[44] = |(datain[135:132] ^ 0);
  assign w133[45] = |(datain[131:128] ^ 15);
  assign w133[46] = |(datain[127:124] ^ 8);
  assign w133[47] = |(datain[123:120] ^ 0);
  assign w133[48] = |(datain[119:116] ^ 15);
  assign w133[49] = |(datain[115:112] ^ 12);
  assign w133[50] = |(datain[111:108] ^ 6);
  assign w133[51] = |(datain[107:104] ^ 4);
  assign w133[52] = |(datain[103:100] ^ 12);
  assign w133[53] = |(datain[99:96] ^ 3);
  assign w133[54] = |(datain[95:92] ^ 8);
  assign w133[55] = |(datain[91:88] ^ 13);
  assign w133[56] = |(datain[87:84] ^ 9);
  assign w133[57] = |(datain[83:80] ^ 6);
  assign w133[58] = |(datain[79:76] ^ 14);
  assign w133[59] = |(datain[75:72] ^ 14);
  assign w133[60] = |(datain[71:68] ^ 0);
  assign w133[61] = |(datain[67:64] ^ 6);
  assign w133[62] = |(datain[63:60] ^ 1);
  assign w133[63] = |(datain[59:56] ^ 14);
  assign w133[64] = |(datain[55:52] ^ 0);
  assign w133[65] = |(datain[51:48] ^ 14);
  assign w133[66] = |(datain[47:44] ^ 1);
  assign w133[67] = |(datain[43:40] ^ 15);
  assign w133[68] = |(datain[39:36] ^ 11);
  assign w133[69] = |(datain[35:32] ^ 4);
  assign w133[70] = |(datain[31:28] ^ 3);
  assign w133[71] = |(datain[27:24] ^ 12);
  assign w133[72] = |(datain[23:20] ^ 11);
  assign w133[73] = |(datain[19:16] ^ 9);
  assign w133[74] = |(datain[15:12] ^ 0);
  assign w133[75] = |(datain[11:8] ^ 3);
  assign comp[133] = ~(|w133);
  wire [74-1:0] w134;
  assign w134[0] = |(datain[311:308] ^ 2);
  assign w134[1] = |(datain[307:304] ^ 1);
  assign w134[2] = |(datain[303:300] ^ 10);
  assign w134[3] = |(datain[299:296] ^ 1);
  assign w134[4] = |(datain[295:292] ^ 7);
  assign w134[5] = |(datain[291:288] ^ 11);
  assign w134[6] = |(datain[287:284] ^ 0);
  assign w134[7] = |(datain[283:280] ^ 7);
  assign w134[8] = |(datain[279:276] ^ 14);
  assign w134[9] = |(datain[275:272] ^ 8);
  assign w134[10] = |(datain[271:268] ^ 3);
  assign w134[11] = |(datain[267:264] ^ 14);
  assign w134[12] = |(datain[263:260] ^ 0);
  assign w134[13] = |(datain[259:256] ^ 0);
  assign w134[14] = |(datain[255:252] ^ 11);
  assign w134[15] = |(datain[251:248] ^ 10);
  assign w134[16] = |(datain[247:244] ^ 8);
  assign w134[17] = |(datain[243:240] ^ 3);
  assign w134[18] = |(datain[239:236] ^ 0);
  assign w134[19] = |(datain[235:232] ^ 7);
  assign w134[20] = |(datain[231:228] ^ 11);
  assign w134[21] = |(datain[227:224] ^ 9);
  assign w134[22] = |(datain[223:220] ^ 1);
  assign w134[23] = |(datain[219:216] ^ 12);
  assign w134[24] = |(datain[215:212] ^ 0);
  assign w134[25] = |(datain[211:208] ^ 0);
  assign w134[26] = |(datain[207:204] ^ 11);
  assign w134[27] = |(datain[203:200] ^ 4);
  assign w134[28] = |(datain[199:196] ^ 4);
  assign w134[29] = |(datain[195:192] ^ 0);
  assign w134[30] = |(datain[191:188] ^ 12);
  assign w134[31] = |(datain[187:184] ^ 13);
  assign w134[32] = |(datain[183:180] ^ 2);
  assign w134[33] = |(datain[179:176] ^ 1);
  assign w134[34] = |(datain[175:172] ^ 2);
  assign w134[35] = |(datain[171:168] ^ 6);
  assign w134[36] = |(datain[167:164] ^ 12);
  assign w134[37] = |(datain[163:160] ^ 7);
  assign w134[38] = |(datain[159:156] ^ 4);
  assign w134[39] = |(datain[155:152] ^ 5);
  assign w134[40] = |(datain[151:148] ^ 1);
  assign w134[41] = |(datain[147:144] ^ 5);
  assign w134[42] = |(datain[143:140] ^ 0);
  assign w134[43] = |(datain[139:136] ^ 0);
  assign w134[44] = |(datain[135:132] ^ 0);
  assign w134[45] = |(datain[131:128] ^ 0);
  assign w134[46] = |(datain[127:124] ^ 2);
  assign w134[47] = |(datain[123:120] ^ 6);
  assign w134[48] = |(datain[119:116] ^ 12);
  assign w134[49] = |(datain[115:112] ^ 7);
  assign w134[50] = |(datain[111:108] ^ 4);
  assign w134[51] = |(datain[107:104] ^ 5);
  assign w134[52] = |(datain[103:100] ^ 1);
  assign w134[53] = |(datain[99:96] ^ 7);
  assign w134[54] = |(datain[95:92] ^ 0);
  assign w134[55] = |(datain[91:88] ^ 0);
  assign w134[56] = |(datain[87:84] ^ 0);
  assign w134[57] = |(datain[83:80] ^ 0);
  assign w134[58] = |(datain[79:76] ^ 11);
  assign w134[59] = |(datain[75:72] ^ 10);
  assign w134[60] = |(datain[71:68] ^ 6);
  assign w134[61] = |(datain[67:64] ^ 7);
  assign w134[62] = |(datain[63:60] ^ 0);
  assign w134[63] = |(datain[59:56] ^ 7);
  assign w134[64] = |(datain[55:52] ^ 11);
  assign w134[65] = |(datain[51:48] ^ 4);
  assign w134[66] = |(datain[47:44] ^ 4);
  assign w134[67] = |(datain[43:40] ^ 0);
  assign w134[68] = |(datain[39:36] ^ 12);
  assign w134[69] = |(datain[35:32] ^ 13);
  assign w134[70] = |(datain[31:28] ^ 2);
  assign w134[71] = |(datain[27:24] ^ 1);
  assign w134[72] = |(datain[23:20] ^ 2);
  assign w134[73] = |(datain[19:16] ^ 6);
  assign comp[134] = ~(|w134);
  wire [76-1:0] w135;
  assign w135[0] = |(datain[311:308] ^ 12);
  assign w135[1] = |(datain[307:304] ^ 7);
  assign w135[2] = |(datain[303:300] ^ 4);
  assign w135[3] = |(datain[299:296] ^ 5);
  assign w135[4] = |(datain[295:292] ^ 1);
  assign w135[5] = |(datain[291:288] ^ 5);
  assign w135[6] = |(datain[287:284] ^ 0);
  assign w135[7] = |(datain[283:280] ^ 0);
  assign w135[8] = |(datain[279:276] ^ 0);
  assign w135[9] = |(datain[275:272] ^ 0);
  assign w135[10] = |(datain[271:268] ^ 2);
  assign w135[11] = |(datain[267:264] ^ 6);
  assign w135[12] = |(datain[263:260] ^ 12);
  assign w135[13] = |(datain[259:256] ^ 7);
  assign w135[14] = |(datain[255:252] ^ 4);
  assign w135[15] = |(datain[251:248] ^ 5);
  assign w135[16] = |(datain[247:244] ^ 1);
  assign w135[17] = |(datain[243:240] ^ 7);
  assign w135[18] = |(datain[239:236] ^ 0);
  assign w135[19] = |(datain[235:232] ^ 0);
  assign w135[20] = |(datain[231:228] ^ 0);
  assign w135[21] = |(datain[227:224] ^ 0);
  assign w135[22] = |(datain[223:220] ^ 11);
  assign w135[23] = |(datain[219:216] ^ 10);
  assign w135[24] = |(datain[215:212] ^ 6);
  assign w135[25] = |(datain[211:208] ^ 7);
  assign w135[26] = |(datain[207:204] ^ 0);
  assign w135[27] = |(datain[203:200] ^ 7);
  assign w135[28] = |(datain[199:196] ^ 11);
  assign w135[29] = |(datain[195:192] ^ 4);
  assign w135[30] = |(datain[191:188] ^ 4);
  assign w135[31] = |(datain[187:184] ^ 0);
  assign w135[32] = |(datain[183:180] ^ 12);
  assign w135[33] = |(datain[179:176] ^ 13);
  assign w135[34] = |(datain[175:172] ^ 2);
  assign w135[35] = |(datain[171:168] ^ 1);
  assign w135[36] = |(datain[167:164] ^ 2);
  assign w135[37] = |(datain[163:160] ^ 6);
  assign w135[38] = |(datain[159:156] ^ 8);
  assign w135[39] = |(datain[155:152] ^ 11);
  assign w135[40] = |(datain[151:148] ^ 4);
  assign w135[41] = |(datain[147:144] ^ 13);
  assign w135[42] = |(datain[143:140] ^ 0);
  assign w135[43] = |(datain[139:136] ^ 13);
  assign w135[44] = |(datain[135:132] ^ 2);
  assign w135[45] = |(datain[131:128] ^ 6);
  assign w135[46] = |(datain[127:124] ^ 8);
  assign w135[47] = |(datain[123:120] ^ 11);
  assign w135[48] = |(datain[119:116] ^ 5);
  assign w135[49] = |(datain[115:112] ^ 5);
  assign w135[50] = |(datain[111:108] ^ 0);
  assign w135[51] = |(datain[107:104] ^ 15);
  assign w135[52] = |(datain[103:100] ^ 13);
  assign w135[53] = |(datain[99:96] ^ 0);
  assign w135[54] = |(datain[95:92] ^ 12);
  assign w135[55] = |(datain[91:88] ^ 14);
  assign w135[56] = |(datain[87:84] ^ 8);
  assign w135[57] = |(datain[83:80] ^ 0);
  assign w135[58] = |(datain[79:76] ^ 12);
  assign w135[59] = |(datain[75:72] ^ 6);
  assign w135[60] = |(datain[71:68] ^ 6);
  assign w135[61] = |(datain[67:64] ^ 4);
  assign w135[62] = |(datain[63:60] ^ 13);
  assign w135[63] = |(datain[59:56] ^ 0);
  assign w135[64] = |(datain[55:52] ^ 12);
  assign w135[65] = |(datain[51:48] ^ 6);
  assign w135[66] = |(datain[47:44] ^ 11);
  assign w135[67] = |(datain[43:40] ^ 8);
  assign w135[68] = |(datain[39:36] ^ 0);
  assign w135[69] = |(datain[35:32] ^ 1);
  assign w135[70] = |(datain[31:28] ^ 5);
  assign w135[71] = |(datain[27:24] ^ 7);
  assign w135[72] = |(datain[23:20] ^ 12);
  assign w135[73] = |(datain[19:16] ^ 13);
  assign w135[74] = |(datain[15:12] ^ 2);
  assign w135[75] = |(datain[11:8] ^ 1);
  assign comp[135] = ~(|w135);
  wire [44-1:0] w136;
  assign w136[0] = |(datain[311:308] ^ 8);
  assign w136[1] = |(datain[307:304] ^ 14);
  assign w136[2] = |(datain[303:300] ^ 13);
  assign w136[3] = |(datain[299:296] ^ 8);
  assign w136[4] = |(datain[295:292] ^ 11);
  assign w136[5] = |(datain[291:288] ^ 14);
  assign w136[6] = |(datain[287:284] ^ 0);
  assign w136[7] = |(datain[283:280] ^ 0);
  assign w136[8] = |(datain[279:276] ^ 0);
  assign w136[9] = |(datain[275:272] ^ 0);
  assign w136[10] = |(datain[271:268] ^ 11);
  assign w136[11] = |(datain[267:264] ^ 0);
  assign w136[12] = |(datain[263:260] ^ 2);
  assign w136[13] = |(datain[259:256] ^ 14);
  assign w136[14] = |(datain[255:252] ^ 11);
  assign w136[15] = |(datain[251:248] ^ 4);
  assign w136[16] = |(datain[247:244] ^ 8);
  assign w136[17] = |(datain[243:240] ^ 0);
  assign w136[18] = |(datain[239:236] ^ 3);
  assign w136[19] = |(datain[235:232] ^ 10);
  assign w136[20] = |(datain[231:228] ^ 0);
  assign w136[21] = |(datain[227:224] ^ 4);
  assign w136[22] = |(datain[223:220] ^ 7);
  assign w136[23] = |(datain[219:216] ^ 5);
  assign w136[24] = |(datain[215:212] ^ 1);
  assign w136[25] = |(datain[211:208] ^ 11);
  assign w136[26] = |(datain[207:204] ^ 11);
  assign w136[27] = |(datain[203:200] ^ 0);
  assign w136[28] = |(datain[199:196] ^ 3);
  assign w136[29] = |(datain[195:192] ^ 10);
  assign w136[30] = |(datain[191:188] ^ 3);
  assign w136[31] = |(datain[187:184] ^ 10);
  assign w136[32] = |(datain[183:180] ^ 4);
  assign w136[33] = |(datain[179:176] ^ 4);
  assign w136[34] = |(datain[175:172] ^ 0);
  assign w136[35] = |(datain[171:168] ^ 1);
  assign w136[36] = |(datain[167:164] ^ 7);
  assign w136[37] = |(datain[163:160] ^ 5);
  assign w136[38] = |(datain[159:156] ^ 1);
  assign w136[39] = |(datain[155:152] ^ 4);
  assign w136[40] = |(datain[151:148] ^ 11);
  assign w136[41] = |(datain[147:144] ^ 0);
  assign w136[42] = |(datain[143:140] ^ 2);
  assign w136[43] = |(datain[139:136] ^ 6);
  assign comp[136] = ~(|w136);
  wire [30-1:0] w137;
  assign w137[0] = |(datain[311:308] ^ 12);
  assign w137[1] = |(datain[307:304] ^ 13);
  assign w137[2] = |(datain[303:300] ^ 2);
  assign w137[3] = |(datain[299:296] ^ 1);
  assign w137[4] = |(datain[295:292] ^ 11);
  assign w137[5] = |(datain[291:288] ^ 9);
  assign w137[6] = |(datain[287:284] ^ 0);
  assign w137[7] = |(datain[283:280] ^ 0);
  assign w137[8] = |(datain[279:276] ^ 12);
  assign w137[9] = |(datain[275:272] ^ 8);
  assign w137[10] = |(datain[271:268] ^ 11);
  assign w137[11] = |(datain[267:264] ^ 11);
  assign w137[12] = |(datain[263:260] ^ 5);
  assign w137[13] = |(datain[259:256] ^ 13);
  assign w137[14] = |(datain[255:252] ^ 2);
  assign w137[15] = |(datain[251:248] ^ 1);
  assign w137[16] = |(datain[247:244] ^ 8);
  assign w137[17] = |(datain[243:240] ^ 9);
  assign w137[18] = |(datain[239:236] ^ 1);
  assign w137[19] = |(datain[235:232] ^ 14);
  assign w137[20] = |(datain[231:228] ^ 4);
  assign w137[21] = |(datain[227:224] ^ 12);
  assign w137[22] = |(datain[223:220] ^ 0);
  assign w137[23] = |(datain[219:216] ^ 0);
  assign w137[24] = |(datain[215:212] ^ 8);
  assign w137[25] = |(datain[211:208] ^ 9);
  assign w137[26] = |(datain[207:204] ^ 0);
  assign w137[27] = |(datain[203:200] ^ 14);
  assign w137[28] = |(datain[199:196] ^ 4);
  assign w137[29] = |(datain[195:192] ^ 14);
  assign comp[137] = ~(|w137);
  wire [74-1:0] w138;
  assign w138[0] = |(datain[311:308] ^ 11);
  assign w138[1] = |(datain[307:304] ^ 8);
  assign w138[2] = |(datain[303:300] ^ 0);
  assign w138[3] = |(datain[299:296] ^ 0);
  assign w138[4] = |(datain[295:292] ^ 4);
  assign w138[5] = |(datain[291:288] ^ 2);
  assign w138[6] = |(datain[287:284] ^ 14);
  assign w138[7] = |(datain[283:280] ^ 8);
  assign w138[8] = |(datain[279:276] ^ 13);
  assign w138[9] = |(datain[275:272] ^ 9);
  assign w138[10] = |(datain[271:268] ^ 15);
  assign w138[11] = |(datain[267:264] ^ 15);
  assign w138[12] = |(datain[263:260] ^ 11);
  assign w138[13] = |(datain[259:256] ^ 4);
  assign w138[14] = |(datain[255:252] ^ 4);
  assign w138[15] = |(datain[251:248] ^ 0);
  assign w138[16] = |(datain[247:244] ^ 8);
  assign w138[17] = |(datain[243:240] ^ 13);
  assign w138[18] = |(datain[239:236] ^ 9);
  assign w138[19] = |(datain[235:232] ^ 6);
  assign w138[20] = |(datain[231:228] ^ 13);
  assign w138[21] = |(datain[227:224] ^ 8);
  assign w138[22] = |(datain[223:220] ^ 0);
  assign w138[23] = |(datain[219:216] ^ 1);
  assign w138[24] = |(datain[215:212] ^ 11);
  assign w138[25] = |(datain[211:208] ^ 9);
  assign w138[26] = |(datain[207:204] ^ 0);
  assign w138[27] = |(datain[203:200] ^ 4);
  assign w138[28] = |(datain[199:196] ^ 0);
  assign w138[29] = |(datain[195:192] ^ 0);
  assign w138[30] = |(datain[191:188] ^ 12);
  assign w138[31] = |(datain[187:184] ^ 13);
  assign w138[32] = |(datain[183:180] ^ 2);
  assign w138[33] = |(datain[179:176] ^ 1);
  assign w138[34] = |(datain[175:172] ^ 14);
  assign w138[35] = |(datain[171:168] ^ 8);
  assign w138[36] = |(datain[167:164] ^ 0);
  assign w138[37] = |(datain[163:160] ^ 14);
  assign w138[38] = |(datain[159:156] ^ 0);
  assign w138[39] = |(datain[155:152] ^ 0);
  assign w138[40] = |(datain[151:148] ^ 11);
  assign w138[41] = |(datain[147:144] ^ 4);
  assign w138[42] = |(datain[143:140] ^ 1);
  assign w138[43] = |(datain[139:136] ^ 10);
  assign w138[44] = |(datain[135:132] ^ 11);
  assign w138[45] = |(datain[131:128] ^ 10);
  assign w138[46] = |(datain[127:124] ^ 8);
  assign w138[47] = |(datain[123:120] ^ 0);
  assign w138[48] = |(datain[119:116] ^ 0);
  assign w138[49] = |(datain[115:112] ^ 0);
  assign w138[50] = |(datain[111:108] ^ 12);
  assign w138[51] = |(datain[107:104] ^ 13);
  assign w138[52] = |(datain[103:100] ^ 2);
  assign w138[53] = |(datain[99:96] ^ 1);
  assign w138[54] = |(datain[95:92] ^ 5);
  assign w138[55] = |(datain[91:88] ^ 8);
  assign w138[56] = |(datain[87:84] ^ 11);
  assign w138[57] = |(datain[83:80] ^ 11);
  assign w138[58] = |(datain[79:76] ^ 0);
  assign w138[59] = |(datain[75:72] ^ 0);
  assign w138[60] = |(datain[71:68] ^ 0);
  assign w138[61] = |(datain[67:64] ^ 1);
  assign w138[62] = |(datain[63:60] ^ 0);
  assign w138[63] = |(datain[59:56] ^ 14);
  assign w138[64] = |(datain[55:52] ^ 5);
  assign w138[65] = |(datain[51:48] ^ 3);
  assign w138[66] = |(datain[47:44] ^ 12);
  assign w138[67] = |(datain[43:40] ^ 11);
  assign w138[68] = |(datain[39:36] ^ 5);
  assign w138[69] = |(datain[35:32] ^ 14);
  assign w138[70] = |(datain[31:28] ^ 5);
  assign w138[71] = |(datain[27:24] ^ 10);
  assign w138[72] = |(datain[23:20] ^ 5);
  assign w138[73] = |(datain[19:16] ^ 9);
  assign comp[138] = ~(|w138);
  wire [74-1:0] w139;
  assign w139[0] = |(datain[311:308] ^ 9);
  assign w139[1] = |(datain[307:304] ^ 6);
  assign w139[2] = |(datain[303:300] ^ 2);
  assign w139[3] = |(datain[299:296] ^ 6);
  assign w139[4] = |(datain[295:292] ^ 0);
  assign w139[5] = |(datain[291:288] ^ 2);
  assign w139[6] = |(datain[287:284] ^ 14);
  assign w139[7] = |(datain[283:280] ^ 8);
  assign w139[8] = |(datain[279:276] ^ 2);
  assign w139[9] = |(datain[275:272] ^ 10);
  assign w139[10] = |(datain[271:268] ^ 0);
  assign w139[11] = |(datain[267:264] ^ 0);
  assign w139[12] = |(datain[263:260] ^ 11);
  assign w139[13] = |(datain[259:256] ^ 4);
  assign w139[14] = |(datain[255:252] ^ 4);
  assign w139[15] = |(datain[251:248] ^ 0);
  assign w139[16] = |(datain[247:244] ^ 11);
  assign w139[17] = |(datain[243:240] ^ 9);
  assign w139[18] = |(datain[239:236] ^ 2);
  assign w139[19] = |(datain[235:232] ^ 10);
  assign w139[20] = |(datain[231:228] ^ 0);
  assign w139[21] = |(datain[227:224] ^ 1);
  assign w139[22] = |(datain[223:220] ^ 8);
  assign w139[23] = |(datain[219:216] ^ 13);
  assign w139[24] = |(datain[215:212] ^ 9);
  assign w139[25] = |(datain[211:208] ^ 6);
  assign w139[26] = |(datain[207:204] ^ 0);
  assign w139[27] = |(datain[203:200] ^ 5);
  assign w139[28] = |(datain[199:196] ^ 0);
  assign w139[29] = |(datain[195:192] ^ 1);
  assign w139[30] = |(datain[191:188] ^ 12);
  assign w139[31] = |(datain[187:184] ^ 13);
  assign w139[32] = |(datain[183:180] ^ 2);
  assign w139[33] = |(datain[179:176] ^ 1);
  assign w139[34] = |(datain[175:172] ^ 14);
  assign w139[35] = |(datain[171:168] ^ 8);
  assign w139[36] = |(datain[167:164] ^ 1);
  assign w139[37] = |(datain[163:160] ^ 12);
  assign w139[38] = |(datain[159:156] ^ 0);
  assign w139[39] = |(datain[155:152] ^ 0);
  assign w139[40] = |(datain[151:148] ^ 11);
  assign w139[41] = |(datain[147:144] ^ 8);
  assign w139[42] = |(datain[143:140] ^ 0);
  assign w139[43] = |(datain[139:136] ^ 0);
  assign w139[44] = |(datain[135:132] ^ 4);
  assign w139[45] = |(datain[131:128] ^ 2);
  assign w139[46] = |(datain[127:124] ^ 2);
  assign w139[47] = |(datain[123:120] ^ 11);
  assign w139[48] = |(datain[119:116] ^ 12);
  assign w139[49] = |(datain[115:112] ^ 9);
  assign w139[50] = |(datain[111:108] ^ 9);
  assign w139[51] = |(datain[107:104] ^ 9);
  assign w139[52] = |(datain[103:100] ^ 12);
  assign w139[53] = |(datain[99:96] ^ 13);
  assign w139[54] = |(datain[95:92] ^ 2);
  assign w139[55] = |(datain[91:88] ^ 1);
  assign w139[56] = |(datain[87:84] ^ 11);
  assign w139[57] = |(datain[83:80] ^ 4);
  assign w139[58] = |(datain[79:76] ^ 4);
  assign w139[59] = |(datain[75:72] ^ 0);
  assign w139[60] = |(datain[71:68] ^ 11);
  assign w139[61] = |(datain[67:64] ^ 9);
  assign w139[62] = |(datain[63:60] ^ 0);
  assign w139[63] = |(datain[59:56] ^ 4);
  assign w139[64] = |(datain[55:52] ^ 0);
  assign w139[65] = |(datain[51:48] ^ 0);
  assign w139[66] = |(datain[47:44] ^ 8);
  assign w139[67] = |(datain[43:40] ^ 13);
  assign w139[68] = |(datain[39:36] ^ 9);
  assign w139[69] = |(datain[35:32] ^ 6);
  assign w139[70] = |(datain[31:28] ^ 11);
  assign w139[71] = |(datain[27:24] ^ 3);
  assign w139[72] = |(datain[23:20] ^ 0);
  assign w139[73] = |(datain[19:16] ^ 1);
  assign comp[139] = ~(|w139);
  wire [76-1:0] w140;
  assign w140[0] = |(datain[311:308] ^ 2);
  assign w140[1] = |(datain[307:304] ^ 13);
  assign w140[2] = |(datain[303:300] ^ 0);
  assign w140[3] = |(datain[299:296] ^ 3);
  assign w140[4] = |(datain[295:292] ^ 0);
  assign w140[5] = |(datain[291:288] ^ 0);
  assign w140[6] = |(datain[287:284] ^ 8);
  assign w140[7] = |(datain[283:280] ^ 9);
  assign w140[8] = |(datain[279:276] ^ 8);
  assign w140[9] = |(datain[275:272] ^ 6);
  assign w140[10] = |(datain[271:268] ^ 11);
  assign w140[11] = |(datain[267:264] ^ 5);
  assign w140[12] = |(datain[263:260] ^ 0);
  assign w140[13] = |(datain[259:256] ^ 1);
  assign w140[14] = |(datain[255:252] ^ 11);
  assign w140[15] = |(datain[251:248] ^ 4);
  assign w140[16] = |(datain[247:244] ^ 4);
  assign w140[17] = |(datain[243:240] ^ 0);
  assign w140[18] = |(datain[239:236] ^ 11);
  assign w140[19] = |(datain[235:232] ^ 9);
  assign w140[20] = |(datain[231:228] ^ 0);
  assign w140[21] = |(datain[227:224] ^ 12);
  assign w140[22] = |(datain[223:220] ^ 0);
  assign w140[23] = |(datain[219:216] ^ 1);
  assign w140[24] = |(datain[215:212] ^ 8);
  assign w140[25] = |(datain[211:208] ^ 13);
  assign w140[26] = |(datain[207:204] ^ 9);
  assign w140[27] = |(datain[203:200] ^ 6);
  assign w140[28] = |(datain[199:196] ^ 0);
  assign w140[29] = |(datain[195:192] ^ 5);
  assign w140[30] = |(datain[191:188] ^ 0);
  assign w140[31] = |(datain[187:184] ^ 1);
  assign w140[32] = |(datain[183:180] ^ 12);
  assign w140[33] = |(datain[179:176] ^ 13);
  assign w140[34] = |(datain[175:172] ^ 2);
  assign w140[35] = |(datain[171:168] ^ 1);
  assign w140[36] = |(datain[167:164] ^ 11);
  assign w140[37] = |(datain[163:160] ^ 8);
  assign w140[38] = |(datain[159:156] ^ 0);
  assign w140[39] = |(datain[155:152] ^ 0);
  assign w140[40] = |(datain[151:148] ^ 4);
  assign w140[41] = |(datain[147:144] ^ 2);
  assign w140[42] = |(datain[143:140] ^ 2);
  assign w140[43] = |(datain[139:136] ^ 11);
  assign w140[44] = |(datain[135:132] ^ 12);
  assign w140[45] = |(datain[131:128] ^ 9);
  assign w140[46] = |(datain[127:124] ^ 9);
  assign w140[47] = |(datain[123:120] ^ 9);
  assign w140[48] = |(datain[119:116] ^ 12);
  assign w140[49] = |(datain[115:112] ^ 13);
  assign w140[50] = |(datain[111:108] ^ 2);
  assign w140[51] = |(datain[107:104] ^ 1);
  assign w140[52] = |(datain[103:100] ^ 11);
  assign w140[53] = |(datain[99:96] ^ 4);
  assign w140[54] = |(datain[95:92] ^ 4);
  assign w140[55] = |(datain[91:88] ^ 0);
  assign w140[56] = |(datain[87:84] ^ 11);
  assign w140[57] = |(datain[83:80] ^ 9);
  assign w140[58] = |(datain[79:76] ^ 0);
  assign w140[59] = |(datain[75:72] ^ 4);
  assign w140[60] = |(datain[71:68] ^ 0);
  assign w140[61] = |(datain[67:64] ^ 0);
  assign w140[62] = |(datain[63:60] ^ 8);
  assign w140[63] = |(datain[59:56] ^ 13);
  assign w140[64] = |(datain[55:52] ^ 9);
  assign w140[65] = |(datain[51:48] ^ 6);
  assign w140[66] = |(datain[47:44] ^ 11);
  assign w140[67] = |(datain[43:40] ^ 4);
  assign w140[68] = |(datain[39:36] ^ 0);
  assign w140[69] = |(datain[35:32] ^ 1);
  assign w140[70] = |(datain[31:28] ^ 12);
  assign w140[71] = |(datain[27:24] ^ 13);
  assign w140[72] = |(datain[23:20] ^ 2);
  assign w140[73] = |(datain[19:16] ^ 1);
  assign w140[74] = |(datain[15:12] ^ 15);
  assign w140[75] = |(datain[11:8] ^ 14);
  assign comp[140] = ~(|w140);
  wire [44-1:0] w141;
  assign w141[0] = |(datain[311:308] ^ 0);
  assign w141[1] = |(datain[307:304] ^ 1);
  assign w141[2] = |(datain[303:300] ^ 4);
  assign w141[3] = |(datain[299:296] ^ 4);
  assign w141[4] = |(datain[295:292] ^ 2);
  assign w141[5] = |(datain[291:288] ^ 5);
  assign w141[6] = |(datain[287:284] ^ 0);
  assign w141[7] = |(datain[283:280] ^ 1);
  assign w141[8] = |(datain[279:276] ^ 4);
  assign w141[9] = |(datain[275:272] ^ 4);
  assign w141[10] = |(datain[271:268] ^ 2);
  assign w141[11] = |(datain[267:264] ^ 7);
  assign w141[12] = |(datain[263:260] ^ 8);
  assign w141[13] = |(datain[259:256] ^ 0);
  assign w141[14] = |(datain[255:252] ^ 3);
  assign w141[15] = |(datain[251:248] ^ 12);
  assign w141[16] = |(datain[247:244] ^ 0);
  assign w141[17] = |(datain[243:240] ^ 0);
  assign w141[18] = |(datain[239:236] ^ 7);
  assign w141[19] = |(datain[235:232] ^ 5);
  assign w141[20] = |(datain[231:228] ^ 0);
  assign w141[21] = |(datain[227:224] ^ 12);
  assign w141[22] = |(datain[223:220] ^ 8);
  assign w141[23] = |(datain[219:216] ^ 11);
  assign w141[24] = |(datain[215:212] ^ 4);
  assign w141[25] = |(datain[211:208] ^ 4);
  assign w141[26] = |(datain[207:204] ^ 0);
  assign w141[27] = |(datain[203:200] ^ 1);
  assign w141[28] = |(datain[199:196] ^ 10);
  assign w141[29] = |(datain[195:192] ^ 3);
  assign w141[30] = |(datain[191:188] ^ 0);
  assign w141[31] = |(datain[187:184] ^ 0);
  assign w141[32] = |(datain[183:180] ^ 0);
  assign w141[33] = |(datain[179:176] ^ 1);
  assign w141[34] = |(datain[175:172] ^ 8);
  assign w141[35] = |(datain[171:168] ^ 10);
  assign w141[36] = |(datain[167:164] ^ 4);
  assign w141[37] = |(datain[163:160] ^ 4);
  assign w141[38] = |(datain[159:156] ^ 0);
  assign w141[39] = |(datain[155:152] ^ 3);
  assign w141[40] = |(datain[151:148] ^ 10);
  assign w141[41] = |(datain[147:144] ^ 2);
  assign w141[42] = |(datain[143:140] ^ 0);
  assign w141[43] = |(datain[139:136] ^ 2);
  assign comp[141] = ~(|w141);
  wire [44-1:0] w142;
  assign w142[0] = |(datain[311:308] ^ 0);
  assign w142[1] = |(datain[307:304] ^ 2);
  assign w142[2] = |(datain[303:300] ^ 11);
  assign w142[3] = |(datain[299:296] ^ 15);
  assign w142[4] = |(datain[295:292] ^ 3);
  assign w142[5] = |(datain[291:288] ^ 4);
  assign w142[6] = |(datain[287:284] ^ 1);
  assign w142[7] = |(datain[283:280] ^ 2);
  assign w142[8] = |(datain[279:276] ^ 12);
  assign w142[9] = |(datain[275:272] ^ 13);
  assign w142[10] = |(datain[271:268] ^ 1);
  assign w142[11] = |(datain[267:264] ^ 3);
  assign w142[12] = |(datain[263:260] ^ 8);
  assign w142[13] = |(datain[259:256] ^ 1);
  assign w142[14] = |(datain[255:252] ^ 15);
  assign w142[15] = |(datain[251:248] ^ 15);
  assign w142[16] = |(datain[247:244] ^ 2);
  assign w142[17] = |(datain[243:240] ^ 1);
  assign w142[18] = |(datain[239:236] ^ 4);
  assign w142[19] = |(datain[235:232] ^ 3);
  assign w142[20] = |(datain[231:228] ^ 7);
  assign w142[21] = |(datain[227:224] ^ 5);
  assign w142[22] = |(datain[223:220] ^ 0);
  assign w142[23] = |(datain[219:216] ^ 3);
  assign w142[24] = |(datain[215:212] ^ 14);
  assign w142[25] = |(datain[211:208] ^ 9);
  assign w142[26] = |(datain[207:204] ^ 2);
  assign w142[27] = |(datain[203:200] ^ 6);
  assign w142[28] = |(datain[199:196] ^ 0);
  assign w142[29] = |(datain[195:192] ^ 1);
  assign w142[30] = |(datain[191:188] ^ 11);
  assign w142[31] = |(datain[187:184] ^ 8);
  assign w142[32] = |(datain[183:180] ^ 2);
  assign w142[33] = |(datain[179:176] ^ 1);
  assign w142[34] = |(datain[175:172] ^ 3);
  assign w142[35] = |(datain[171:168] ^ 5);
  assign w142[36] = |(datain[167:164] ^ 12);
  assign w142[37] = |(datain[163:160] ^ 13);
  assign w142[38] = |(datain[159:156] ^ 2);
  assign w142[39] = |(datain[155:152] ^ 1);
  assign w142[40] = |(datain[151:148] ^ 8);
  assign w142[41] = |(datain[147:144] ^ 9);
  assign w142[42] = |(datain[143:140] ^ 1);
  assign w142[43] = |(datain[139:136] ^ 14);
  assign comp[142] = ~(|w142);
  wire [56-1:0] w143;
  assign w143[0] = |(datain[311:308] ^ 9);
  assign w143[1] = |(datain[307:304] ^ 6);
  assign w143[2] = |(datain[303:300] ^ 8);
  assign w143[3] = |(datain[299:296] ^ 5);
  assign w143[4] = |(datain[295:292] ^ 0);
  assign w143[5] = |(datain[291:288] ^ 5);
  assign w143[6] = |(datain[287:284] ^ 8);
  assign w143[7] = |(datain[283:280] ^ 13);
  assign w143[8] = |(datain[279:276] ^ 11);
  assign w143[9] = |(datain[275:272] ^ 6);
  assign w143[10] = |(datain[271:268] ^ 1);
  assign w143[11] = |(datain[267:264] ^ 12);
  assign w143[12] = |(datain[263:260] ^ 0);
  assign w143[13] = |(datain[259:256] ^ 0);
  assign w143[14] = |(datain[255:252] ^ 11);
  assign w143[15] = |(datain[251:248] ^ 9);
  assign w143[16] = |(datain[247:244] ^ 11);
  assign w143[17] = |(datain[243:240] ^ 2);
  assign w143[18] = |(datain[239:236] ^ 0);
  assign w143[19] = |(datain[235:232] ^ 2);
  assign w143[20] = |(datain[231:228] ^ 3);
  assign w143[21] = |(datain[227:224] ^ 1);
  assign w143[22] = |(datain[223:220] ^ 1);
  assign w143[23] = |(datain[219:216] ^ 4);
  assign w143[24] = |(datain[215:212] ^ 4);
  assign w143[25] = |(datain[211:208] ^ 6);
  assign w143[26] = |(datain[207:204] ^ 4);
  assign w143[27] = |(datain[203:200] ^ 6);
  assign w143[28] = |(datain[199:196] ^ 14);
  assign w143[29] = |(datain[195:192] ^ 2);
  assign w143[30] = |(datain[191:188] ^ 15);
  assign w143[31] = |(datain[187:184] ^ 10);
  assign w143[32] = |(datain[183:180] ^ 12);
  assign w143[33] = |(datain[179:176] ^ 3);
  assign w143[34] = |(datain[175:172] ^ 14);
  assign w143[35] = |(datain[171:168] ^ 8);
  assign w143[36] = |(datain[167:164] ^ 0);
  assign w143[37] = |(datain[163:160] ^ 0);
  assign w143[38] = |(datain[159:156] ^ 0);
  assign w143[39] = |(datain[155:152] ^ 0);
  assign w143[40] = |(datain[151:148] ^ 5);
  assign w143[41] = |(datain[147:144] ^ 13);
  assign w143[42] = |(datain[143:140] ^ 8);
  assign w143[43] = |(datain[139:136] ^ 1);
  assign w143[44] = |(datain[135:132] ^ 14);
  assign w143[45] = |(datain[131:128] ^ 13);
  assign w143[46] = |(datain[127:124] ^ 11);
  assign w143[47] = |(datain[123:120] ^ 14);
  assign w143[48] = |(datain[119:116] ^ 0);
  assign w143[49] = |(datain[115:112] ^ 5);
  assign w143[50] = |(datain[111:108] ^ 14);
  assign w143[51] = |(datain[107:104] ^ 11);
  assign w143[52] = |(datain[103:100] ^ 0);
  assign w143[53] = |(datain[99:96] ^ 0);
  assign w143[54] = |(datain[95:92] ^ 12);
  assign w143[55] = |(datain[91:88] ^ 3);
  assign comp[143] = ~(|w143);
  wire [76-1:0] w144;
  assign w144[0] = |(datain[311:308] ^ 2);
  assign w144[1] = |(datain[307:304] ^ 6);
  assign w144[2] = |(datain[303:300] ^ 8);
  assign w144[3] = |(datain[299:296] ^ 9);
  assign w144[4] = |(datain[295:292] ^ 4);
  assign w144[5] = |(datain[291:288] ^ 5);
  assign w144[6] = |(datain[287:284] ^ 1);
  assign w144[7] = |(datain[283:280] ^ 5);
  assign w144[8] = |(datain[279:276] ^ 11);
  assign w144[9] = |(datain[275:272] ^ 4);
  assign w144[10] = |(datain[271:268] ^ 4);
  assign w144[11] = |(datain[267:264] ^ 0);
  assign w144[12] = |(datain[263:260] ^ 11);
  assign w144[13] = |(datain[259:256] ^ 9);
  assign w144[14] = |(datain[255:252] ^ 10);
  assign w144[15] = |(datain[251:248] ^ 7);
  assign w144[16] = |(datain[247:244] ^ 0);
  assign w144[17] = |(datain[243:240] ^ 1);
  assign w144[18] = |(datain[239:236] ^ 11);
  assign w144[19] = |(datain[235:232] ^ 10);
  assign w144[20] = |(datain[231:228] ^ 10);
  assign w144[21] = |(datain[227:224] ^ 11);
  assign w144[22] = |(datain[223:220] ^ 0);
  assign w144[23] = |(datain[219:216] ^ 2);
  assign w144[24] = |(datain[215:212] ^ 9);
  assign w144[25] = |(datain[211:208] ^ 12);
  assign w144[26] = |(datain[207:204] ^ 2);
  assign w144[27] = |(datain[203:200] ^ 14);
  assign w144[28] = |(datain[199:196] ^ 15);
  assign w144[29] = |(datain[195:192] ^ 15);
  assign w144[30] = |(datain[191:188] ^ 1);
  assign w144[31] = |(datain[187:184] ^ 14);
  assign w144[32] = |(datain[183:180] ^ 9);
  assign w144[33] = |(datain[179:176] ^ 13);
  assign w144[34] = |(datain[175:172] ^ 0);
  assign w144[35] = |(datain[171:168] ^ 2);
  assign w144[36] = |(datain[167:164] ^ 3);
  assign w144[37] = |(datain[163:160] ^ 3);
  assign w144[38] = |(datain[159:156] ^ 12);
  assign w144[39] = |(datain[155:152] ^ 0);
  assign w144[40] = |(datain[151:148] ^ 2);
  assign w144[41] = |(datain[147:144] ^ 6);
  assign w144[42] = |(datain[143:140] ^ 8);
  assign w144[43] = |(datain[139:136] ^ 9);
  assign w144[44] = |(datain[135:132] ^ 4);
  assign w144[45] = |(datain[131:128] ^ 5);
  assign w144[46] = |(datain[127:124] ^ 1);
  assign w144[47] = |(datain[123:120] ^ 5);
  assign w144[48] = |(datain[119:116] ^ 11);
  assign w144[49] = |(datain[115:112] ^ 4);
  assign w144[50] = |(datain[111:108] ^ 4);
  assign w144[51] = |(datain[107:104] ^ 0);
  assign w144[52] = |(datain[103:100] ^ 11);
  assign w144[53] = |(datain[99:96] ^ 9);
  assign w144[54] = |(datain[95:92] ^ 0);
  assign w144[55] = |(datain[91:88] ^ 3);
  assign w144[56] = |(datain[87:84] ^ 0);
  assign w144[57] = |(datain[83:80] ^ 0);
  assign w144[58] = |(datain[79:76] ^ 2);
  assign w144[59] = |(datain[75:72] ^ 9);
  assign w144[60] = |(datain[71:68] ^ 0);
  assign w144[61] = |(datain[67:64] ^ 14);
  assign w144[62] = |(datain[63:60] ^ 10);
  assign w144[63] = |(datain[59:56] ^ 2);
  assign w144[64] = |(datain[55:52] ^ 0);
  assign w144[65] = |(datain[51:48] ^ 2);
  assign w144[66] = |(datain[47:44] ^ 11);
  assign w144[67] = |(datain[43:40] ^ 10);
  assign w144[68] = |(datain[39:36] ^ 10);
  assign w144[69] = |(datain[35:32] ^ 1);
  assign w144[70] = |(datain[31:28] ^ 0);
  assign w144[71] = |(datain[27:24] ^ 2);
  assign w144[72] = |(datain[23:20] ^ 9);
  assign w144[73] = |(datain[19:16] ^ 12);
  assign w144[74] = |(datain[15:12] ^ 2);
  assign w144[75] = |(datain[11:8] ^ 14);
  assign comp[144] = ~(|w144);
  wire [76-1:0] w145;
  assign w145[0] = |(datain[311:308] ^ 4);
  assign w145[1] = |(datain[307:304] ^ 9);
  assign w145[2] = |(datain[303:300] ^ 0);
  assign w145[3] = |(datain[299:296] ^ 1);
  assign w145[4] = |(datain[295:292] ^ 5);
  assign w145[5] = |(datain[291:288] ^ 9);
  assign w145[6] = |(datain[287:284] ^ 5);
  assign w145[7] = |(datain[283:280] ^ 8);
  assign w145[8] = |(datain[279:276] ^ 11);
  assign w145[9] = |(datain[275:272] ^ 4);
  assign w145[10] = |(datain[271:268] ^ 4);
  assign w145[11] = |(datain[267:264] ^ 0);
  assign w145[12] = |(datain[263:260] ^ 11);
  assign w145[13] = |(datain[259:256] ^ 9);
  assign w145[14] = |(datain[255:252] ^ 1);
  assign w145[15] = |(datain[251:248] ^ 3);
  assign w145[16] = |(datain[247:244] ^ 0);
  assign w145[17] = |(datain[243:240] ^ 3);
  assign w145[18] = |(datain[239:236] ^ 11);
  assign w145[19] = |(datain[235:232] ^ 10);
  assign w145[20] = |(datain[231:228] ^ 0);
  assign w145[21] = |(datain[227:224] ^ 0);
  assign w145[22] = |(datain[223:220] ^ 0);
  assign w145[23] = |(datain[219:216] ^ 1);
  assign w145[24] = |(datain[215:212] ^ 9);
  assign w145[25] = |(datain[211:208] ^ 12);
  assign w145[26] = |(datain[207:204] ^ 2);
  assign w145[27] = |(datain[203:200] ^ 14);
  assign w145[28] = |(datain[199:196] ^ 15);
  assign w145[29] = |(datain[195:192] ^ 15);
  assign w145[30] = |(datain[191:188] ^ 1);
  assign w145[31] = |(datain[187:184] ^ 14);
  assign w145[32] = |(datain[183:180] ^ 1);
  assign w145[33] = |(datain[179:176] ^ 9);
  assign w145[34] = |(datain[175:172] ^ 0);
  assign w145[35] = |(datain[171:168] ^ 1);
  assign w145[36] = |(datain[167:164] ^ 7);
  assign w145[37] = |(datain[163:160] ^ 2);
  assign w145[38] = |(datain[159:156] ^ 1);
  assign w145[39] = |(datain[155:152] ^ 13);
  assign w145[40] = |(datain[151:148] ^ 11);
  assign w145[41] = |(datain[147:144] ^ 8);
  assign w145[42] = |(datain[143:140] ^ 0);
  assign w145[43] = |(datain[139:136] ^ 0);
  assign w145[44] = |(datain[135:132] ^ 4);
  assign w145[45] = |(datain[131:128] ^ 2);
  assign w145[46] = |(datain[127:124] ^ 3);
  assign w145[47] = |(datain[123:120] ^ 3);
  assign w145[48] = |(datain[119:116] ^ 12);
  assign w145[49] = |(datain[115:112] ^ 9);
  assign w145[50] = |(datain[111:108] ^ 3);
  assign w145[51] = |(datain[107:104] ^ 3);
  assign w145[52] = |(datain[103:100] ^ 13);
  assign w145[53] = |(datain[99:96] ^ 2);
  assign w145[54] = |(datain[95:92] ^ 9);
  assign w145[55] = |(datain[91:88] ^ 12);
  assign w145[56] = |(datain[87:84] ^ 2);
  assign w145[57] = |(datain[83:80] ^ 14);
  assign w145[58] = |(datain[79:76] ^ 15);
  assign w145[59] = |(datain[75:72] ^ 15);
  assign w145[60] = |(datain[71:68] ^ 1);
  assign w145[61] = |(datain[67:64] ^ 14);
  assign w145[62] = |(datain[63:60] ^ 1);
  assign w145[63] = |(datain[59:56] ^ 9);
  assign w145[64] = |(datain[55:52] ^ 0);
  assign w145[65] = |(datain[51:48] ^ 1);
  assign w145[66] = |(datain[47:44] ^ 7);
  assign w145[67] = |(datain[43:40] ^ 2);
  assign w145[68] = |(datain[39:36] ^ 0);
  assign w145[69] = |(datain[35:32] ^ 14);
  assign w145[70] = |(datain[31:28] ^ 11);
  assign w145[71] = |(datain[27:24] ^ 10);
  assign w145[72] = |(datain[23:20] ^ 1);
  assign w145[73] = |(datain[19:16] ^ 13);
  assign w145[74] = |(datain[15:12] ^ 0);
  assign w145[75] = |(datain[11:8] ^ 1);
  assign comp[145] = ~(|w145);
  wire [76-1:0] w146;
  assign w146[0] = |(datain[311:308] ^ 1);
  assign w146[1] = |(datain[307:304] ^ 9);
  assign w146[2] = |(datain[303:300] ^ 0);
  assign w146[3] = |(datain[299:296] ^ 1);
  assign w146[4] = |(datain[295:292] ^ 7);
  assign w146[5] = |(datain[291:288] ^ 2);
  assign w146[6] = |(datain[287:284] ^ 0);
  assign w146[7] = |(datain[283:280] ^ 14);
  assign w146[8] = |(datain[279:276] ^ 11);
  assign w146[9] = |(datain[275:272] ^ 10);
  assign w146[10] = |(datain[271:268] ^ 1);
  assign w146[11] = |(datain[267:264] ^ 13);
  assign w146[12] = |(datain[263:260] ^ 0);
  assign w146[13] = |(datain[259:256] ^ 1);
  assign w146[14] = |(datain[255:252] ^ 11);
  assign w146[15] = |(datain[251:248] ^ 9);
  assign w146[16] = |(datain[247:244] ^ 2);
  assign w146[17] = |(datain[243:240] ^ 0);
  assign w146[18] = |(datain[239:236] ^ 0);
  assign w146[19] = |(datain[235:232] ^ 0);
  assign w146[20] = |(datain[231:228] ^ 11);
  assign w146[21] = |(datain[227:224] ^ 4);
  assign w146[22] = |(datain[223:220] ^ 4);
  assign w146[23] = |(datain[219:216] ^ 0);
  assign w146[24] = |(datain[215:212] ^ 9);
  assign w146[25] = |(datain[211:208] ^ 12);
  assign w146[26] = |(datain[207:204] ^ 2);
  assign w146[27] = |(datain[203:200] ^ 14);
  assign w146[28] = |(datain[199:196] ^ 15);
  assign w146[29] = |(datain[195:192] ^ 15);
  assign w146[30] = |(datain[191:188] ^ 1);
  assign w146[31] = |(datain[187:184] ^ 14);
  assign w146[32] = |(datain[183:180] ^ 1);
  assign w146[33] = |(datain[179:176] ^ 9);
  assign w146[34] = |(datain[175:172] ^ 0);
  assign w146[35] = |(datain[171:168] ^ 1);
  assign w146[36] = |(datain[167:164] ^ 2);
  assign w146[37] = |(datain[163:160] ^ 14);
  assign w146[38] = |(datain[159:156] ^ 8);
  assign w146[39] = |(datain[155:152] ^ 11);
  assign w146[40] = |(datain[151:148] ^ 0);
  assign w146[41] = |(datain[147:144] ^ 14);
  assign w146[42] = |(datain[143:140] ^ 4);
  assign w146[43] = |(datain[139:136] ^ 5);
  assign w146[44] = |(datain[135:132] ^ 0);
  assign w146[45] = |(datain[131:128] ^ 1);
  assign w146[46] = |(datain[127:124] ^ 2);
  assign w146[47] = |(datain[123:120] ^ 14);
  assign w146[48] = |(datain[119:116] ^ 8);
  assign w146[49] = |(datain[115:112] ^ 11);
  assign w146[50] = |(datain[111:108] ^ 1);
  assign w146[51] = |(datain[107:104] ^ 6);
  assign w146[52] = |(datain[103:100] ^ 4);
  assign w146[53] = |(datain[99:96] ^ 7);
  assign w146[54] = |(datain[95:92] ^ 0);
  assign w146[55] = |(datain[91:88] ^ 1);
  assign w146[56] = |(datain[87:84] ^ 11);
  assign w146[57] = |(datain[83:80] ^ 8);
  assign w146[58] = |(datain[79:76] ^ 0);
  assign w146[59] = |(datain[75:72] ^ 1);
  assign w146[60] = |(datain[71:68] ^ 5);
  assign w146[61] = |(datain[67:64] ^ 7);
  assign w146[62] = |(datain[63:60] ^ 9);
  assign w146[63] = |(datain[59:56] ^ 12);
  assign w146[64] = |(datain[55:52] ^ 2);
  assign w146[65] = |(datain[51:48] ^ 14);
  assign w146[66] = |(datain[47:44] ^ 15);
  assign w146[67] = |(datain[43:40] ^ 15);
  assign w146[68] = |(datain[39:36] ^ 1);
  assign w146[69] = |(datain[35:32] ^ 14);
  assign w146[70] = |(datain[31:28] ^ 1);
  assign w146[71] = |(datain[27:24] ^ 9);
  assign w146[72] = |(datain[23:20] ^ 0);
  assign w146[73] = |(datain[19:16] ^ 1);
  assign w146[74] = |(datain[15:12] ^ 11);
  assign w146[75] = |(datain[11:8] ^ 4);
  assign comp[146] = ~(|w146);
  wire [74-1:0] w147;
  assign w147[0] = |(datain[311:308] ^ 11);
  assign w147[1] = |(datain[307:304] ^ 4);
  assign w147[2] = |(datain[303:300] ^ 6);
  assign w147[3] = |(datain[299:296] ^ 6);
  assign w147[4] = |(datain[295:292] ^ 12);
  assign w147[5] = |(datain[291:288] ^ 15);
  assign w147[6] = |(datain[287:284] ^ 5);
  assign w147[7] = |(datain[283:280] ^ 10);
  assign w147[8] = |(datain[279:276] ^ 1);
  assign w147[9] = |(datain[275:272] ^ 15);
  assign w147[10] = |(datain[271:268] ^ 14);
  assign w147[11] = |(datain[267:264] ^ 11);
  assign w147[12] = |(datain[263:260] ^ 15);
  assign w147[13] = |(datain[259:256] ^ 6);
  assign w147[14] = |(datain[255:252] ^ 11);
  assign w147[15] = |(datain[251:248] ^ 10);
  assign w147[16] = |(datain[247:244] ^ 8);
  assign w147[17] = |(datain[243:240] ^ 0);
  assign w147[18] = |(datain[239:236] ^ 0);
  assign w147[19] = |(datain[235:232] ^ 0);
  assign w147[20] = |(datain[231:228] ^ 12);
  assign w147[21] = |(datain[227:224] ^ 13);
  assign w147[22] = |(datain[223:220] ^ 6);
  assign w147[23] = |(datain[219:216] ^ 6);
  assign w147[24] = |(datain[215:212] ^ 12);
  assign w147[25] = |(datain[211:208] ^ 3);
  assign w147[26] = |(datain[207:204] ^ 11);
  assign w147[27] = |(datain[203:200] ^ 4);
  assign w147[28] = |(datain[199:196] ^ 4);
  assign w147[29] = |(datain[195:192] ^ 0);
  assign w147[30] = |(datain[191:188] ^ 12);
  assign w147[31] = |(datain[187:184] ^ 13);
  assign w147[32] = |(datain[183:180] ^ 2);
  assign w147[33] = |(datain[179:176] ^ 1);
  assign w147[34] = |(datain[175:172] ^ 12);
  assign w147[35] = |(datain[171:168] ^ 3);
  assign w147[36] = |(datain[167:164] ^ 14);
  assign w147[37] = |(datain[163:160] ^ 8);
  assign w147[38] = |(datain[159:156] ^ 6);
  assign w147[39] = |(datain[155:152] ^ 11);
  assign w147[40] = |(datain[151:148] ^ 0);
  assign w147[41] = |(datain[147:144] ^ 1);
  assign w147[42] = |(datain[143:140] ^ 11);
  assign w147[43] = |(datain[139:136] ^ 10);
  assign w147[44] = |(datain[135:132] ^ 0);
  assign w147[45] = |(datain[131:128] ^ 0);
  assign w147[46] = |(datain[127:124] ^ 0);
  assign w147[47] = |(datain[123:120] ^ 6);
  assign w147[48] = |(datain[119:116] ^ 11);
  assign w147[49] = |(datain[115:112] ^ 9);
  assign w147[50] = |(datain[111:108] ^ 0);
  assign w147[51] = |(datain[107:104] ^ 0);
  assign w147[52] = |(datain[103:100] ^ 0);
  assign w147[53] = |(datain[99:96] ^ 6);
  assign w147[54] = |(datain[95:92] ^ 14);
  assign w147[55] = |(datain[91:88] ^ 8);
  assign w147[56] = |(datain[87:84] ^ 14);
  assign w147[57] = |(datain[83:80] ^ 15);
  assign w147[58] = |(datain[79:76] ^ 15);
  assign w147[59] = |(datain[75:72] ^ 15);
  assign w147[60] = |(datain[71:68] ^ 12);
  assign w147[61] = |(datain[67:64] ^ 3);
  assign w147[62] = |(datain[63:60] ^ 11);
  assign w147[63] = |(datain[59:56] ^ 4);
  assign w147[64] = |(datain[55:52] ^ 4);
  assign w147[65] = |(datain[51:48] ^ 2);
  assign w147[66] = |(datain[47:44] ^ 2);
  assign w147[67] = |(datain[43:40] ^ 11);
  assign w147[68] = |(datain[39:36] ^ 12);
  assign w147[69] = |(datain[35:32] ^ 9);
  assign w147[70] = |(datain[31:28] ^ 2);
  assign w147[71] = |(datain[27:24] ^ 11);
  assign w147[72] = |(datain[23:20] ^ 13);
  assign w147[73] = |(datain[19:16] ^ 2);
  assign comp[147] = ~(|w147);
  wire [34-1:0] w148;
  assign w148[0] = |(datain[311:308] ^ 15);
  assign w148[1] = |(datain[307:304] ^ 15);
  assign w148[2] = |(datain[303:300] ^ 15);
  assign w148[3] = |(datain[299:296] ^ 15);
  assign w148[4] = |(datain[295:292] ^ 7);
  assign w148[5] = |(datain[291:288] ^ 2);
  assign w148[6] = |(datain[287:284] ^ 0);
  assign w148[7] = |(datain[283:280] ^ 3);
  assign w148[8] = |(datain[279:276] ^ 10);
  assign w148[9] = |(datain[275:272] ^ 3);
  assign w148[10] = |(datain[271:268] ^ 9);
  assign w148[11] = |(datain[267:264] ^ 11);
  assign w148[12] = |(datain[263:260] ^ 0);
  assign w148[13] = |(datain[259:256] ^ 0);
  assign w148[14] = |(datain[255:252] ^ 10);
  assign w148[15] = |(datain[251:248] ^ 1);
  assign w148[16] = |(datain[247:244] ^ 9);
  assign w148[17] = |(datain[243:240] ^ 11);
  assign w148[18] = |(datain[239:236] ^ 0);
  assign w148[19] = |(datain[235:232] ^ 0);
  assign w148[20] = |(datain[231:228] ^ 3);
  assign w148[21] = |(datain[227:224] ^ 13);
  assign w148[22] = |(datain[223:220] ^ 15);
  assign w148[23] = |(datain[219:216] ^ 15);
  assign w148[24] = |(datain[215:212] ^ 15);
  assign w148[25] = |(datain[211:208] ^ 15);
  assign w148[26] = |(datain[207:204] ^ 7);
  assign w148[27] = |(datain[203:200] ^ 4);
  assign w148[28] = |(datain[199:196] ^ 1);
  assign w148[29] = |(datain[195:192] ^ 15);
  assign w148[30] = |(datain[191:188] ^ 11);
  assign w148[31] = |(datain[187:184] ^ 0);
  assign w148[32] = |(datain[183:180] ^ 0);
  assign w148[33] = |(datain[179:176] ^ 0);
  assign comp[148] = ~(|w148);
  wire [30-1:0] w149;
  assign w149[0] = |(datain[311:308] ^ 14);
  assign w149[1] = |(datain[307:304] ^ 1);
  assign w149[2] = |(datain[303:300] ^ 15);
  assign w149[3] = |(datain[299:296] ^ 15);
  assign w149[4] = |(datain[295:292] ^ 14);
  assign w149[5] = |(datain[291:288] ^ 8);
  assign w149[6] = |(datain[287:284] ^ 13);
  assign w149[7] = |(datain[283:280] ^ 1);
  assign w149[8] = |(datain[279:276] ^ 15);
  assign w149[9] = |(datain[275:272] ^ 15);
  assign w149[10] = |(datain[271:268] ^ 0);
  assign w149[11] = |(datain[267:264] ^ 7);
  assign w149[12] = |(datain[263:260] ^ 9);
  assign w149[13] = |(datain[259:256] ^ 12);
  assign w149[14] = |(datain[255:252] ^ 3);
  assign w149[15] = |(datain[251:248] ^ 3);
  assign w149[16] = |(datain[247:244] ^ 12);
  assign w149[17] = |(datain[243:240] ^ 0);
  assign w149[18] = |(datain[239:236] ^ 8);
  assign w149[19] = |(datain[235:232] ^ 14);
  assign w149[20] = |(datain[231:228] ^ 12);
  assign w149[21] = |(datain[227:224] ^ 0);
  assign w149[22] = |(datain[223:220] ^ 2);
  assign w149[23] = |(datain[219:216] ^ 6);
  assign w149[24] = |(datain[215:212] ^ 15);
  assign w149[25] = |(datain[211:208] ^ 15);
  assign w149[26] = |(datain[207:204] ^ 1);
  assign w149[27] = |(datain[203:200] ^ 14);
  assign w149[28] = |(datain[199:196] ^ 0);
  assign w149[29] = |(datain[195:192] ^ 4);
  assign comp[149] = ~(|w149);
  wire [28-1:0] w150;
  assign w150[0] = |(datain[311:308] ^ 14);
  assign w150[1] = |(datain[307:304] ^ 8);
  assign w150[2] = |(datain[303:300] ^ 13);
  assign w150[3] = |(datain[299:296] ^ 1);
  assign w150[4] = |(datain[295:292] ^ 15);
  assign w150[5] = |(datain[291:288] ^ 15);
  assign w150[6] = |(datain[287:284] ^ 0);
  assign w150[7] = |(datain[283:280] ^ 7);
  assign w150[8] = |(datain[279:276] ^ 9);
  assign w150[9] = |(datain[275:272] ^ 12);
  assign w150[10] = |(datain[271:268] ^ 3);
  assign w150[11] = |(datain[267:264] ^ 3);
  assign w150[12] = |(datain[263:260] ^ 12);
  assign w150[13] = |(datain[259:256] ^ 0);
  assign w150[14] = |(datain[255:252] ^ 8);
  assign w150[15] = |(datain[251:248] ^ 14);
  assign w150[16] = |(datain[247:244] ^ 12);
  assign w150[17] = |(datain[243:240] ^ 0);
  assign w150[18] = |(datain[239:236] ^ 2);
  assign w150[19] = |(datain[235:232] ^ 6);
  assign w150[20] = |(datain[231:228] ^ 15);
  assign w150[21] = |(datain[227:224] ^ 15);
  assign w150[22] = |(datain[223:220] ^ 1);
  assign w150[23] = |(datain[219:216] ^ 14);
  assign w150[24] = |(datain[215:212] ^ 0);
  assign w150[25] = |(datain[211:208] ^ 4);
  assign w150[26] = |(datain[207:204] ^ 0);
  assign w150[27] = |(datain[203:200] ^ 0);
  assign comp[150] = ~(|w150);
  wire [28-1:0] w151;
  assign w151[0] = |(datain[311:308] ^ 14);
  assign w151[1] = |(datain[307:304] ^ 12);
  assign w151[2] = |(datain[303:300] ^ 11);
  assign w151[3] = |(datain[299:296] ^ 14);
  assign w151[4] = |(datain[295:292] ^ 3);
  assign w151[5] = |(datain[291:288] ^ 12);
  assign w151[6] = |(datain[287:284] ^ 0);
  assign w151[7] = |(datain[283:280] ^ 1);
  assign w151[8] = |(datain[279:276] ^ 11);
  assign w151[9] = |(datain[275:272] ^ 15);
  assign w151[10] = |(datain[271:268] ^ 0);
  assign w151[11] = |(datain[267:264] ^ 0);
  assign w151[12] = |(datain[263:260] ^ 0);
  assign w151[13] = |(datain[259:256] ^ 0);
  assign w151[14] = |(datain[255:252] ^ 11);
  assign w151[15] = |(datain[251:248] ^ 9);
  assign w151[16] = |(datain[247:244] ^ 1);
  assign w151[17] = |(datain[243:240] ^ 0);
  assign w151[18] = |(datain[239:236] ^ 0);
  assign w151[19] = |(datain[235:232] ^ 0);
  assign w151[20] = |(datain[231:228] ^ 15);
  assign w151[21] = |(datain[227:224] ^ 12);
  assign w151[22] = |(datain[223:220] ^ 15);
  assign w151[23] = |(datain[219:216] ^ 2);
  assign w151[24] = |(datain[215:212] ^ 10);
  assign w151[25] = |(datain[211:208] ^ 4);
  assign w151[26] = |(datain[207:204] ^ 14);
  assign w151[27] = |(datain[203:200] ^ 9);
  assign comp[151] = ~(|w151);
  wire [26-1:0] w152;
  assign w152[0] = |(datain[311:308] ^ 12);
  assign w152[1] = |(datain[307:304] ^ 0);
  assign w152[2] = |(datain[303:300] ^ 12);
  assign w152[3] = |(datain[299:296] ^ 11);
  assign w152[4] = |(datain[295:292] ^ 11);
  assign w152[5] = |(datain[291:288] ^ 14);
  assign w152[6] = |(datain[287:284] ^ 0);
  assign w152[7] = |(datain[283:280] ^ 6);
  assign w152[8] = |(datain[279:276] ^ 0);
  assign w152[9] = |(datain[275:272] ^ 0);
  assign w152[10] = |(datain[271:268] ^ 10);
  assign w152[11] = |(datain[267:264] ^ 13);
  assign w152[12] = |(datain[263:260] ^ 3);
  assign w152[13] = |(datain[259:256] ^ 13);
  assign w152[14] = |(datain[255:252] ^ 9);
  assign w152[15] = |(datain[251:248] ^ 2);
  assign w152[16] = |(datain[247:244] ^ 0);
  assign w152[17] = |(datain[243:240] ^ 1);
  assign w152[18] = |(datain[239:236] ^ 7);
  assign w152[19] = |(datain[235:232] ^ 4);
  assign w152[20] = |(datain[231:228] ^ 13);
  assign w152[21] = |(datain[227:224] ^ 13);
  assign w152[22] = |(datain[223:220] ^ 3);
  assign w152[23] = |(datain[219:216] ^ 13);
  assign w152[24] = |(datain[215:212] ^ 7);
  assign w152[25] = |(datain[211:208] ^ 9);
  assign comp[152] = ~(|w152);
  wire [28-1:0] w153;
  assign w153[0] = |(datain[311:308] ^ 0);
  assign w153[1] = |(datain[307:304] ^ 6);
  assign w153[2] = |(datain[303:300] ^ 15);
  assign w153[3] = |(datain[299:296] ^ 0);
  assign w153[4] = |(datain[295:292] ^ 0);
  assign w153[5] = |(datain[291:288] ^ 4);
  assign w153[6] = |(datain[287:284] ^ 15);
  assign w153[7] = |(datain[283:280] ^ 3);
  assign w153[8] = |(datain[279:276] ^ 10);
  assign w153[9] = |(datain[275:272] ^ 4);
  assign w153[10] = |(datain[271:268] ^ 2);
  assign w153[11] = |(datain[267:264] ^ 6);
  assign w153[12] = |(datain[263:260] ^ 12);
  assign w153[13] = |(datain[259:256] ^ 6);
  assign w153[14] = |(datain[255:252] ^ 0);
  assign w153[15] = |(datain[251:248] ^ 6);
  assign w153[16] = |(datain[247:244] ^ 15);
  assign w153[17] = |(datain[243:240] ^ 2);
  assign w153[18] = |(datain[239:236] ^ 0);
  assign w153[19] = |(datain[235:232] ^ 4);
  assign w153[20] = |(datain[231:228] ^ 12);
  assign w153[21] = |(datain[227:224] ^ 11);
  assign w153[22] = |(datain[223:220] ^ 5);
  assign w153[23] = |(datain[219:216] ^ 15);
  assign w153[24] = |(datain[215:212] ^ 0);
  assign w153[25] = |(datain[211:208] ^ 7);
  assign w153[26] = |(datain[207:204] ^ 12);
  assign w153[27] = |(datain[203:200] ^ 3);
  assign comp[153] = ~(|w153);
  wire [28-1:0] w154;
  assign w154[0] = |(datain[311:308] ^ 8);
  assign w154[1] = |(datain[307:304] ^ 13);
  assign w154[2] = |(datain[303:300] ^ 1);
  assign w154[3] = |(datain[299:296] ^ 6);
  assign w154[4] = |(datain[295:292] ^ 5);
  assign w154[5] = |(datain[291:288] ^ 3);
  assign w154[6] = |(datain[287:284] ^ 0);
  assign w154[7] = |(datain[283:280] ^ 1);
  assign w154[8] = |(datain[279:276] ^ 11);
  assign w154[9] = |(datain[275:272] ^ 8);
  assign w154[10] = |(datain[271:268] ^ 2);
  assign w154[11] = |(datain[267:264] ^ 1);
  assign w154[12] = |(datain[263:260] ^ 2);
  assign w154[13] = |(datain[259:256] ^ 5);
  assign w154[14] = |(datain[255:252] ^ 12);
  assign w154[15] = |(datain[251:248] ^ 13);
  assign w154[16] = |(datain[247:244] ^ 2);
  assign w154[17] = |(datain[243:240] ^ 1);
  assign w154[18] = |(datain[239:236] ^ 5);
  assign w154[19] = |(datain[235:232] ^ 10);
  assign w154[20] = |(datain[231:228] ^ 11);
  assign w154[21] = |(datain[227:224] ^ 11);
  assign w154[22] = |(datain[223:220] ^ 11);
  assign w154[23] = |(datain[219:216] ^ 0);
  assign w154[24] = |(datain[215:212] ^ 0);
  assign w154[25] = |(datain[211:208] ^ 2);
  assign w154[26] = |(datain[207:204] ^ 0);
  assign w154[27] = |(datain[203:200] ^ 1);
  assign comp[154] = ~(|w154);
  wire [32-1:0] w155;
  assign w155[0] = |(datain[311:308] ^ 8);
  assign w155[1] = |(datain[307:304] ^ 11);
  assign w155[2] = |(datain[303:300] ^ 3);
  assign w155[3] = |(datain[299:296] ^ 5);
  assign w155[4] = |(datain[295:292] ^ 8);
  assign w155[5] = |(datain[291:288] ^ 9);
  assign w155[6] = |(datain[287:284] ^ 3);
  assign w155[7] = |(datain[283:280] ^ 6);
  assign w155[8] = |(datain[279:276] ^ 0);
  assign w155[9] = |(datain[275:272] ^ 0);
  assign w155[10] = |(datain[271:268] ^ 0);
  assign w155[11] = |(datain[267:264] ^ 1);
  assign w155[12] = |(datain[263:260] ^ 8);
  assign w155[13] = |(datain[259:256] ^ 11);
  assign w155[14] = |(datain[255:252] ^ 7);
  assign w155[15] = |(datain[251:248] ^ 5);
  assign w155[16] = |(datain[247:244] ^ 0);
  assign w155[17] = |(datain[243:240] ^ 2);
  assign w155[18] = |(datain[239:236] ^ 8);
  assign w155[19] = |(datain[235:232] ^ 9);
  assign w155[20] = |(datain[231:228] ^ 3);
  assign w155[21] = |(datain[227:224] ^ 6);
  assign w155[22] = |(datain[223:220] ^ 0);
  assign w155[23] = |(datain[219:216] ^ 2);
  assign w155[24] = |(datain[215:212] ^ 0);
  assign w155[25] = |(datain[211:208] ^ 1);
  assign w155[26] = |(datain[207:204] ^ 12);
  assign w155[27] = |(datain[203:200] ^ 7);
  assign w155[28] = |(datain[199:196] ^ 4);
  assign w155[29] = |(datain[195:192] ^ 5);
  assign w155[30] = |(datain[191:188] ^ 1);
  assign w155[31] = |(datain[187:184] ^ 4);
  assign comp[155] = ~(|w155);
  wire [30-1:0] w156;
  assign w156[0] = |(datain[311:308] ^ 0);
  assign w156[1] = |(datain[307:304] ^ 2);
  assign w156[2] = |(datain[303:300] ^ 12);
  assign w156[3] = |(datain[299:296] ^ 13);
  assign w156[4] = |(datain[295:292] ^ 2);
  assign w156[5] = |(datain[291:288] ^ 1);
  assign w156[6] = |(datain[287:284] ^ 11);
  assign w156[7] = |(datain[283:280] ^ 8);
  assign w156[8] = |(datain[279:276] ^ 1);
  assign w156[9] = |(datain[275:272] ^ 3);
  assign w156[10] = |(datain[271:268] ^ 2);
  assign w156[11] = |(datain[267:264] ^ 5);
  assign w156[12] = |(datain[263:260] ^ 11);
  assign w156[13] = |(datain[259:256] ^ 10);
  assign w156[14] = |(datain[255:252] ^ 14);
  assign w156[15] = |(datain[251:248] ^ 11);
  assign w156[16] = |(datain[247:244] ^ 0);
  assign w156[17] = |(datain[243:240] ^ 1);
  assign w156[18] = |(datain[239:236] ^ 12);
  assign w156[19] = |(datain[235:232] ^ 13);
  assign w156[20] = |(datain[231:228] ^ 2);
  assign w156[21] = |(datain[227:224] ^ 1);
  assign w156[22] = |(datain[223:220] ^ 8);
  assign w156[23] = |(datain[219:216] ^ 14);
  assign w156[24] = |(datain[215:212] ^ 0);
  assign w156[25] = |(datain[211:208] ^ 6);
  assign w156[26] = |(datain[207:204] ^ 2);
  assign w156[27] = |(datain[203:200] ^ 13);
  assign w156[28] = |(datain[199:196] ^ 0);
  assign w156[29] = |(datain[195:192] ^ 0);
  assign comp[156] = ~(|w156);
  wire [32-1:0] w157;
  assign w157[0] = |(datain[311:308] ^ 11);
  assign w157[1] = |(datain[307:304] ^ 15);
  assign w157[2] = |(datain[303:300] ^ 0);
  assign w157[3] = |(datain[299:296] ^ 0);
  assign w157[4] = |(datain[295:292] ^ 0);
  assign w157[5] = |(datain[291:288] ^ 1);
  assign w157[6] = |(datain[287:284] ^ 11);
  assign w157[7] = |(datain[283:280] ^ 14);
  assign w157[8] = |(datain[279:276] ^ 4);
  assign w157[9] = |(datain[275:272] ^ 0);
  assign w157[10] = |(datain[271:268] ^ 0);
  assign w157[11] = |(datain[267:264] ^ 6);
  assign w157[12] = |(datain[263:260] ^ 0);
  assign w157[13] = |(datain[259:256] ^ 3);
  assign w157[14] = |(datain[255:252] ^ 15);
  assign w157[15] = |(datain[251:248] ^ 7);
  assign w157[16] = |(datain[247:244] ^ 2);
  assign w157[17] = |(datain[243:240] ^ 14);
  assign w157[18] = |(datain[239:236] ^ 8);
  assign w157[19] = |(datain[235:232] ^ 11);
  assign w157[20] = |(datain[231:228] ^ 8);
  assign w157[21] = |(datain[227:224] ^ 13);
  assign w157[22] = |(datain[223:220] ^ 0);
  assign w157[23] = |(datain[219:216] ^ 15);
  assign w157[24] = |(datain[215:212] ^ 0);
  assign w157[25] = |(datain[211:208] ^ 0);
  assign w157[26] = |(datain[207:204] ^ 12);
  assign w157[27] = |(datain[203:200] ^ 13);
  assign w157[28] = |(datain[199:196] ^ 2);
  assign w157[29] = |(datain[195:192] ^ 1);
  assign w157[30] = |(datain[191:188] ^ 8);
  assign w157[31] = |(datain[187:184] ^ 12);
  assign comp[157] = ~(|w157);
  wire [76-1:0] w158;
  assign w158[0] = |(datain[311:308] ^ 12);
  assign w158[1] = |(datain[307:304] ^ 0);
  assign w158[2] = |(datain[303:300] ^ 11);
  assign w158[3] = |(datain[299:296] ^ 4);
  assign w158[4] = |(datain[295:292] ^ 4);
  assign w158[5] = |(datain[291:288] ^ 2);
  assign w158[6] = |(datain[287:284] ^ 3);
  assign w158[7] = |(datain[283:280] ^ 3);
  assign w158[8] = |(datain[279:276] ^ 12);
  assign w158[9] = |(datain[275:272] ^ 9);
  assign w158[10] = |(datain[271:268] ^ 9);
  assign w158[11] = |(datain[267:264] ^ 9);
  assign w158[12] = |(datain[263:260] ^ 12);
  assign w158[13] = |(datain[259:256] ^ 13);
  assign w158[14] = |(datain[255:252] ^ 2);
  assign w158[15] = |(datain[251:248] ^ 1);
  assign w158[16] = |(datain[247:244] ^ 11);
  assign w158[17] = |(datain[243:240] ^ 4);
  assign w158[18] = |(datain[239:236] ^ 4);
  assign w158[19] = |(datain[235:232] ^ 0);
  assign w158[20] = |(datain[231:228] ^ 11);
  assign w158[21] = |(datain[227:224] ^ 9);
  assign w158[22] = |(datain[223:220] ^ 1);
  assign w158[23] = |(datain[219:216] ^ 0);
  assign w158[24] = |(datain[215:212] ^ 0);
  assign w158[25] = |(datain[211:208] ^ 1);
  assign w158[26] = |(datain[207:204] ^ 11);
  assign w158[27] = |(datain[203:200] ^ 10);
  assign w158[28] = |(datain[199:196] ^ 0);
  assign w158[29] = |(datain[195:192] ^ 0);
  assign w158[30] = |(datain[191:188] ^ 0);
  assign w158[31] = |(datain[187:184] ^ 1);
  assign w158[32] = |(datain[183:180] ^ 12);
  assign w158[33] = |(datain[179:176] ^ 13);
  assign w158[34] = |(datain[175:172] ^ 2);
  assign w158[35] = |(datain[171:168] ^ 1);
  assign w158[36] = |(datain[167:164] ^ 11);
  assign w158[37] = |(datain[163:160] ^ 4);
  assign w158[38] = |(datain[159:156] ^ 3);
  assign w158[39] = |(datain[155:152] ^ 14);
  assign w158[40] = |(datain[151:148] ^ 12);
  assign w158[41] = |(datain[147:144] ^ 13);
  assign w158[42] = |(datain[143:140] ^ 2);
  assign w158[43] = |(datain[139:136] ^ 1);
  assign w158[44] = |(datain[135:132] ^ 12);
  assign w158[45] = |(datain[131:128] ^ 13);
  assign w158[46] = |(datain[127:124] ^ 2);
  assign w158[47] = |(datain[123:120] ^ 0);
  assign w158[48] = |(datain[119:116] ^ 6);
  assign w158[49] = |(datain[115:112] ^ 13);
  assign w158[50] = |(datain[111:108] ^ 6);
  assign w158[51] = |(datain[107:104] ^ 1);
  assign w158[52] = |(datain[103:100] ^ 6);
  assign w158[53] = |(datain[99:96] ^ 11);
  assign w158[54] = |(datain[95:92] ^ 6);
  assign w158[55] = |(datain[91:88] ^ 9);
  assign w158[56] = |(datain[87:84] ^ 6);
  assign w158[57] = |(datain[83:80] ^ 14);
  assign w158[58] = |(datain[79:76] ^ 6);
  assign w158[59] = |(datain[75:72] ^ 7);
  assign w158[60] = |(datain[71:68] ^ 2);
  assign w158[61] = |(datain[67:64] ^ 0);
  assign w158[62] = |(datain[63:60] ^ 5);
  assign w158[63] = |(datain[59:56] ^ 6);
  assign w158[64] = |(datain[55:52] ^ 6);
  assign w158[65] = |(datain[51:48] ^ 9);
  assign w158[66] = |(datain[47:44] ^ 7);
  assign w158[67] = |(datain[43:40] ^ 2);
  assign w158[68] = |(datain[39:36] ^ 5);
  assign w158[69] = |(datain[35:32] ^ 5);
  assign w158[70] = |(datain[31:28] ^ 4);
  assign w158[71] = |(datain[27:24] ^ 3);
  assign w158[72] = |(datain[23:20] ^ 7);
  assign w158[73] = |(datain[19:16] ^ 4);
  assign w158[74] = |(datain[15:12] ^ 4);
  assign w158[75] = |(datain[11:8] ^ 9);
  assign comp[158] = ~(|w158);
  wire [74-1:0] w159;
  assign w159[0] = |(datain[311:308] ^ 0);
  assign w159[1] = |(datain[307:304] ^ 11);
  assign w159[2] = |(datain[303:300] ^ 11);
  assign w159[3] = |(datain[299:296] ^ 14);
  assign w159[4] = |(datain[295:292] ^ 15);
  assign w159[5] = |(datain[291:288] ^ 7);
  assign w159[6] = |(datain[287:284] ^ 0);
  assign w159[7] = |(datain[283:280] ^ 5);
  assign w159[8] = |(datain[279:276] ^ 11);
  assign w159[9] = |(datain[275:272] ^ 9);
  assign w159[10] = |(datain[271:268] ^ 13);
  assign w159[11] = |(datain[267:264] ^ 8);
  assign w159[12] = |(datain[263:260] ^ 0);
  assign w159[13] = |(datain[259:256] ^ 4);
  assign w159[14] = |(datain[255:252] ^ 11);
  assign w159[15] = |(datain[251:248] ^ 10);
  assign w159[16] = |(datain[247:244] ^ 0);
  assign w159[17] = |(datain[243:240] ^ 3);
  assign w159[18] = |(datain[239:236] ^ 0);
  assign w159[19] = |(datain[235:232] ^ 1);
  assign w159[20] = |(datain[231:228] ^ 14);
  assign w159[21] = |(datain[227:224] ^ 8);
  assign w159[22] = |(datain[223:220] ^ 9);
  assign w159[23] = |(datain[219:216] ^ 5);
  assign w159[24] = |(datain[215:212] ^ 0);
  assign w159[25] = |(datain[211:208] ^ 1);
  assign w159[26] = |(datain[207:204] ^ 11);
  assign w159[27] = |(datain[203:200] ^ 4);
  assign w159[28] = |(datain[199:196] ^ 4);
  assign w159[29] = |(datain[195:192] ^ 0);
  assign w159[30] = |(datain[191:188] ^ 12);
  assign w159[31] = |(datain[187:184] ^ 13);
  assign w159[32] = |(datain[183:180] ^ 2);
  assign w159[33] = |(datain[179:176] ^ 1);
  assign w159[34] = |(datain[175:172] ^ 0);
  assign w159[35] = |(datain[171:168] ^ 7);
  assign w159[36] = |(datain[167:164] ^ 5);
  assign w159[37] = |(datain[163:160] ^ 15);
  assign w159[38] = |(datain[159:156] ^ 11);
  assign w159[39] = |(datain[155:152] ^ 4);
  assign w159[40] = |(datain[151:148] ^ 4);
  assign w159[41] = |(datain[147:144] ^ 0);
  assign w159[42] = |(datain[143:140] ^ 11);
  assign w159[43] = |(datain[139:136] ^ 9);
  assign w159[44] = |(datain[135:132] ^ 1);
  assign w159[45] = |(datain[131:128] ^ 12);
  assign w159[46] = |(datain[127:124] ^ 0);
  assign w159[47] = |(datain[123:120] ^ 0);
  assign w159[48] = |(datain[119:116] ^ 11);
  assign w159[49] = |(datain[115:112] ^ 10);
  assign w159[50] = |(datain[111:108] ^ 13);
  assign w159[51] = |(datain[107:104] ^ 11);
  assign w159[52] = |(datain[103:100] ^ 0);
  assign w159[53] = |(datain[99:96] ^ 5);
  assign w159[54] = |(datain[95:92] ^ 12);
  assign w159[55] = |(datain[91:88] ^ 13);
  assign w159[56] = |(datain[87:84] ^ 2);
  assign w159[57] = |(datain[83:80] ^ 1);
  assign w159[58] = |(datain[79:76] ^ 14);
  assign w159[59] = |(datain[75:72] ^ 8);
  assign w159[60] = |(datain[71:68] ^ 6);
  assign w159[61] = |(datain[67:64] ^ 12);
  assign w159[62] = |(datain[63:60] ^ 0);
  assign w159[63] = |(datain[59:56] ^ 1);
  assign w159[64] = |(datain[55:52] ^ 11);
  assign w159[65] = |(datain[51:48] ^ 4);
  assign w159[66] = |(datain[47:44] ^ 4);
  assign w159[67] = |(datain[43:40] ^ 0);
  assign w159[68] = |(datain[39:36] ^ 11);
  assign w159[69] = |(datain[35:32] ^ 9);
  assign w159[70] = |(datain[31:28] ^ 1);
  assign w159[71] = |(datain[27:24] ^ 10);
  assign w159[72] = |(datain[23:20] ^ 0);
  assign w159[73] = |(datain[19:16] ^ 0);
  assign comp[159] = ~(|w159);
  wire [76-1:0] w160;
  assign w160[0] = |(datain[311:308] ^ 12);
  assign w160[1] = |(datain[307:304] ^ 13);
  assign w160[2] = |(datain[303:300] ^ 2);
  assign w160[3] = |(datain[299:296] ^ 1);
  assign w160[4] = |(datain[295:292] ^ 9);
  assign w160[5] = |(datain[291:288] ^ 3);
  assign w160[6] = |(datain[287:284] ^ 12);
  assign w160[7] = |(datain[283:280] ^ 3);
  assign w160[8] = |(datain[279:276] ^ 11);
  assign w160[9] = |(datain[275:272] ^ 4);
  assign w160[10] = |(datain[271:268] ^ 3);
  assign w160[11] = |(datain[267:264] ^ 14);
  assign w160[12] = |(datain[263:260] ^ 12);
  assign w160[13] = |(datain[259:256] ^ 13);
  assign w160[14] = |(datain[255:252] ^ 2);
  assign w160[15] = |(datain[251:248] ^ 1);
  assign w160[16] = |(datain[247:244] ^ 12);
  assign w160[17] = |(datain[243:240] ^ 3);
  assign w160[18] = |(datain[239:236] ^ 11);
  assign w160[19] = |(datain[235:232] ^ 4);
  assign w160[20] = |(datain[231:228] ^ 3);
  assign w160[21] = |(datain[227:224] ^ 15);
  assign w160[22] = |(datain[223:220] ^ 12);
  assign w160[23] = |(datain[219:216] ^ 13);
  assign w160[24] = |(datain[215:212] ^ 2);
  assign w160[25] = |(datain[211:208] ^ 1);
  assign w160[26] = |(datain[207:204] ^ 12);
  assign w160[27] = |(datain[203:200] ^ 3);
  assign w160[28] = |(datain[199:196] ^ 11);
  assign w160[29] = |(datain[195:192] ^ 4);
  assign w160[30] = |(datain[191:188] ^ 4);
  assign w160[31] = |(datain[187:184] ^ 0);
  assign w160[32] = |(datain[183:180] ^ 12);
  assign w160[33] = |(datain[179:176] ^ 13);
  assign w160[34] = |(datain[175:172] ^ 2);
  assign w160[35] = |(datain[171:168] ^ 1);
  assign w160[36] = |(datain[167:164] ^ 12);
  assign w160[37] = |(datain[163:160] ^ 3);
  assign w160[38] = |(datain[159:156] ^ 11);
  assign w160[39] = |(datain[155:152] ^ 4);
  assign w160[40] = |(datain[151:148] ^ 4);
  assign w160[41] = |(datain[147:144] ^ 3);
  assign w160[42] = |(datain[143:140] ^ 12);
  assign w160[43] = |(datain[139:136] ^ 13);
  assign w160[44] = |(datain[135:132] ^ 2);
  assign w160[45] = |(datain[131:128] ^ 1);
  assign w160[46] = |(datain[127:124] ^ 12);
  assign w160[47] = |(datain[123:120] ^ 3);
  assign w160[48] = |(datain[119:116] ^ 11);
  assign w160[49] = |(datain[115:112] ^ 4);
  assign w160[50] = |(datain[111:108] ^ 5);
  assign w160[51] = |(datain[107:104] ^ 6);
  assign w160[52] = |(datain[103:100] ^ 12);
  assign w160[53] = |(datain[99:96] ^ 13);
  assign w160[54] = |(datain[95:92] ^ 2);
  assign w160[55] = |(datain[91:88] ^ 1);
  assign w160[56] = |(datain[87:84] ^ 12);
  assign w160[57] = |(datain[83:80] ^ 3);
  assign w160[58] = |(datain[79:76] ^ 9);
  assign w160[59] = |(datain[75:72] ^ 12);
  assign w160[60] = |(datain[71:68] ^ 3);
  assign w160[61] = |(datain[67:64] ^ 13);
  assign w160[62] = |(datain[63:60] ^ 10);
  assign w160[63] = |(datain[59:56] ^ 11);
  assign w160[64] = |(datain[55:52] ^ 6);
  assign w160[65] = |(datain[51:48] ^ 3);
  assign w160[66] = |(datain[47:44] ^ 7);
  assign w160[67] = |(datain[43:40] ^ 5);
  assign w160[68] = |(datain[39:36] ^ 0);
  assign w160[69] = |(datain[35:32] ^ 4);
  assign w160[70] = |(datain[31:28] ^ 3);
  assign w160[71] = |(datain[27:24] ^ 3);
  assign w160[72] = |(datain[23:20] ^ 15);
  assign w160[73] = |(datain[19:16] ^ 6);
  assign w160[74] = |(datain[15:12] ^ 9);
  assign w160[75] = |(datain[11:8] ^ 13);
  assign comp[160] = ~(|w160);
  wire [32-1:0] w161;
  assign w161[0] = |(datain[311:308] ^ 5);
  assign w161[1] = |(datain[307:304] ^ 11);
  assign w161[2] = |(datain[303:300] ^ 8);
  assign w161[3] = |(datain[299:296] ^ 1);
  assign w161[4] = |(datain[295:292] ^ 12);
  assign w161[5] = |(datain[291:288] ^ 3);
  assign w161[6] = |(datain[287:284] ^ 1);
  assign w161[7] = |(datain[283:280] ^ 0);
  assign w161[8] = |(datain[279:276] ^ 0);
  assign w161[9] = |(datain[275:272] ^ 0);
  assign w161[10] = |(datain[271:268] ^ 11);
  assign w161[11] = |(datain[267:264] ^ 9);
  assign w161[12] = |(datain[263:260] ^ 7);
  assign w161[13] = |(datain[259:256] ^ 0);
  assign w161[14] = |(datain[255:252] ^ 0);
  assign w161[15] = |(datain[251:248] ^ 6);
  assign w161[16] = |(datain[247:244] ^ 3);
  assign w161[17] = |(datain[243:240] ^ 3);
  assign w161[18] = |(datain[239:236] ^ 15);
  assign w161[19] = |(datain[235:232] ^ 6);
  assign w161[20] = |(datain[231:228] ^ 8);
  assign w161[21] = |(datain[227:224] ^ 0);
  assign w161[22] = |(datain[223:220] ^ 3);
  assign w161[23] = |(datain[219:216] ^ 0);
  assign w161[24] = |(datain[215:212] ^ 11);
  assign w161[25] = |(datain[211:208] ^ 13);
  assign w161[26] = |(datain[207:204] ^ 4);
  assign w161[27] = |(datain[203:200] ^ 6);
  assign w161[28] = |(datain[199:196] ^ 14);
  assign w161[29] = |(datain[195:192] ^ 2);
  assign w161[30] = |(datain[191:188] ^ 15);
  assign w161[31] = |(datain[187:184] ^ 10);
  assign comp[161] = ~(|w161);
  wire [48-1:0] w162;
  assign w162[0] = |(datain[311:308] ^ 7);
  assign w162[1] = |(datain[307:304] ^ 15);
  assign w162[2] = |(datain[303:300] ^ 0);
  assign w162[3] = |(datain[299:296] ^ 8);
  assign w162[4] = |(datain[295:292] ^ 0);
  assign w162[5] = |(datain[291:288] ^ 3);
  assign w162[6] = |(datain[287:284] ^ 7);
  assign w162[7] = |(datain[283:280] ^ 5);
  assign w162[8] = |(datain[279:276] ^ 0);
  assign w162[9] = |(datain[275:272] ^ 8);
  assign w162[10] = |(datain[271:268] ^ 8);
  assign w162[11] = |(datain[267:264] ^ 11);
  assign w162[12] = |(datain[263:260] ^ 13);
  assign w162[13] = |(datain[259:256] ^ 8);
  assign w162[14] = |(datain[255:252] ^ 8);
  assign w162[15] = |(datain[251:248] ^ 3);
  assign w162[16] = |(datain[247:244] ^ 7);
  assign w162[17] = |(datain[243:240] ^ 15);
  assign w162[18] = |(datain[239:236] ^ 0);
  assign w162[19] = |(datain[235:232] ^ 6);
  assign w162[20] = |(datain[231:228] ^ 0);
  assign w162[21] = |(datain[227:224] ^ 1);
  assign w162[22] = |(datain[223:220] ^ 7);
  assign w162[23] = |(datain[219:216] ^ 4);
  assign w162[24] = |(datain[215:212] ^ 0);
  assign w162[25] = |(datain[211:208] ^ 15);
  assign w162[26] = |(datain[207:204] ^ 8);
  assign w162[27] = |(datain[203:200] ^ 11);
  assign w162[28] = |(datain[199:196] ^ 5);
  assign w162[29] = |(datain[195:192] ^ 14);
  assign w162[30] = |(datain[191:188] ^ 15);
  assign w162[31] = |(datain[187:184] ^ 12);
  assign w162[32] = |(datain[183:180] ^ 8);
  assign w162[33] = |(datain[179:176] ^ 3);
  assign w162[34] = |(datain[175:172] ^ 7);
  assign w162[35] = |(datain[171:168] ^ 15);
  assign w162[36] = |(datain[167:164] ^ 0);
  assign w162[37] = |(datain[163:160] ^ 12);
  assign w162[38] = |(datain[159:156] ^ 0);
  assign w162[39] = |(datain[155:152] ^ 5);
  assign w162[40] = |(datain[151:148] ^ 7);
  assign w162[41] = |(datain[147:144] ^ 5);
  assign w162[42] = |(datain[143:140] ^ 4);
  assign w162[43] = |(datain[139:136] ^ 1);
  assign w162[44] = |(datain[135:132] ^ 8);
  assign w162[45] = |(datain[131:128] ^ 3);
  assign w162[46] = |(datain[127:124] ^ 7);
  assign w162[47] = |(datain[123:120] ^ 15);
  assign comp[162] = ~(|w162);
  wire [26-1:0] w163;
  assign w163[0] = |(datain[311:308] ^ 0);
  assign w163[1] = |(datain[307:304] ^ 15);
  assign w163[2] = |(datain[303:300] ^ 8);
  assign w163[3] = |(datain[299:296] ^ 13);
  assign w163[4] = |(datain[295:292] ^ 11);
  assign w163[5] = |(datain[291:288] ^ 7);
  assign w163[6] = |(datain[287:284] ^ 4);
  assign w163[7] = |(datain[283:280] ^ 13);
  assign w163[8] = |(datain[279:276] ^ 0);
  assign w163[9] = |(datain[275:272] ^ 1);
  assign w163[10] = |(datain[271:268] ^ 11);
  assign w163[11] = |(datain[267:264] ^ 12);
  assign w163[12] = |(datain[263:260] ^ 8);
  assign w163[13] = |(datain[259:256] ^ 2);
  assign w163[14] = |(datain[255:252] ^ 0);
  assign w163[15] = |(datain[251:248] ^ 6);
  assign w163[16] = |(datain[247:244] ^ 3);
  assign w163[17] = |(datain[243:240] ^ 1);
  assign w163[18] = |(datain[239:236] ^ 3);
  assign w163[19] = |(datain[235:232] ^ 4);
  assign w163[20] = |(datain[231:228] ^ 3);
  assign w163[21] = |(datain[227:224] ^ 1);
  assign w163[22] = |(datain[223:220] ^ 2);
  assign w163[23] = |(datain[219:216] ^ 4);
  assign w163[24] = |(datain[215:212] ^ 4);
  assign w163[25] = |(datain[211:208] ^ 6);
  assign comp[163] = ~(|w163);
  wire [30-1:0] w164;
  assign w164[0] = |(datain[311:308] ^ 8);
  assign w164[1] = |(datain[307:304] ^ 13);
  assign w164[2] = |(datain[303:300] ^ 11);
  assign w164[3] = |(datain[299:296] ^ 7);
  assign w164[4] = |(datain[295:292] ^ 4);
  assign w164[5] = |(datain[291:288] ^ 11);
  assign w164[6] = |(datain[287:284] ^ 0);
  assign w164[7] = |(datain[283:280] ^ 1);
  assign w164[8] = |(datain[279:276] ^ 11);
  assign w164[9] = |(datain[275:272] ^ 12);
  assign w164[10] = |(datain[271:268] ^ 8);
  assign w164[11] = |(datain[267:264] ^ 8);
  assign w164[12] = |(datain[263:260] ^ 0);
  assign w164[13] = |(datain[259:256] ^ 6);
  assign w164[14] = |(datain[255:252] ^ 3);
  assign w164[15] = |(datain[251:248] ^ 1);
  assign w164[16] = |(datain[247:244] ^ 3);
  assign w164[17] = |(datain[243:240] ^ 4);
  assign w164[18] = |(datain[239:236] ^ 3);
  assign w164[19] = |(datain[235:232] ^ 1);
  assign w164[20] = |(datain[231:228] ^ 2);
  assign w164[21] = |(datain[227:224] ^ 4);
  assign w164[22] = |(datain[223:220] ^ 4);
  assign w164[23] = |(datain[219:216] ^ 6);
  assign w164[24] = |(datain[215:212] ^ 4);
  assign w164[25] = |(datain[211:208] ^ 12);
  assign w164[26] = |(datain[207:204] ^ 7);
  assign w164[27] = |(datain[203:200] ^ 5);
  assign w164[28] = |(datain[199:196] ^ 15);
  assign w164[29] = |(datain[195:192] ^ 8);
  assign comp[164] = ~(|w164);
  wire [76-1:0] w165;
  assign w165[0] = |(datain[311:308] ^ 5);
  assign w165[1] = |(datain[307:304] ^ 9);
  assign w165[2] = |(datain[303:300] ^ 8);
  assign w165[3] = |(datain[299:296] ^ 13);
  assign w165[4] = |(datain[295:292] ^ 9);
  assign w165[5] = |(datain[291:288] ^ 6);
  assign w165[6] = |(datain[287:284] ^ 7);
  assign w165[7] = |(datain[283:280] ^ 15);
  assign w165[8] = |(datain[279:276] ^ 0);
  assign w165[9] = |(datain[275:272] ^ 5);
  assign w165[10] = |(datain[271:268] ^ 12);
  assign w165[11] = |(datain[267:264] ^ 13);
  assign w165[12] = |(datain[263:260] ^ 2);
  assign w165[13] = |(datain[259:256] ^ 1);
  assign w165[14] = |(datain[255:252] ^ 3);
  assign w165[15] = |(datain[251:248] ^ 2);
  assign w165[16] = |(datain[247:244] ^ 12);
  assign w165[17] = |(datain[243:240] ^ 0);
  assign w165[18] = |(datain[239:236] ^ 14);
  assign w165[19] = |(datain[235:232] ^ 8);
  assign w165[20] = |(datain[231:228] ^ 2);
  assign w165[21] = |(datain[227:224] ^ 9);
  assign w165[22] = |(datain[223:220] ^ 0);
  assign w165[23] = |(datain[219:216] ^ 0);
  assign w165[24] = |(datain[215:212] ^ 8);
  assign w165[25] = |(datain[211:208] ^ 13);
  assign w165[26] = |(datain[207:204] ^ 9);
  assign w165[27] = |(datain[203:200] ^ 6);
  assign w165[28] = |(datain[199:196] ^ 13);
  assign w165[29] = |(datain[195:192] ^ 15);
  assign w165[30] = |(datain[191:188] ^ 0);
  assign w165[31] = |(datain[187:184] ^ 4);
  assign w165[32] = |(datain[183:180] ^ 12);
  assign w165[33] = |(datain[179:176] ^ 13);
  assign w165[34] = |(datain[175:172] ^ 2);
  assign w165[35] = |(datain[171:168] ^ 1);
  assign w165[36] = |(datain[167:164] ^ 5);
  assign w165[37] = |(datain[163:160] ^ 10);
  assign w165[38] = |(datain[159:156] ^ 5);
  assign w165[39] = |(datain[155:152] ^ 9);
  assign w165[40] = |(datain[151:148] ^ 8);
  assign w165[41] = |(datain[147:144] ^ 0);
  assign w165[42] = |(datain[143:140] ^ 14);
  assign w165[43] = |(datain[139:136] ^ 1);
  assign w165[44] = |(datain[135:132] ^ 14);
  assign w165[45] = |(datain[131:128] ^ 0);
  assign w165[46] = |(datain[127:124] ^ 8);
  assign w165[47] = |(datain[123:120] ^ 0);
  assign w165[48] = |(datain[119:116] ^ 12);
  assign w165[49] = |(datain[115:112] ^ 9);
  assign w165[50] = |(datain[111:108] ^ 1);
  assign w165[51] = |(datain[107:104] ^ 13);
  assign w165[52] = |(datain[103:100] ^ 11);
  assign w165[53] = |(datain[99:96] ^ 8);
  assign w165[54] = |(datain[95:92] ^ 0);
  assign w165[55] = |(datain[91:88] ^ 1);
  assign w165[56] = |(datain[87:84] ^ 5);
  assign w165[57] = |(datain[83:80] ^ 7);
  assign w165[58] = |(datain[79:76] ^ 12);
  assign w165[59] = |(datain[75:72] ^ 13);
  assign w165[60] = |(datain[71:68] ^ 2);
  assign w165[61] = |(datain[67:64] ^ 1);
  assign w165[62] = |(datain[63:60] ^ 1);
  assign w165[63] = |(datain[59:56] ^ 15);
  assign w165[64] = |(datain[55:52] ^ 5);
  assign w165[65] = |(datain[51:48] ^ 10);
  assign w165[66] = |(datain[47:44] ^ 5);
  assign w165[67] = |(datain[43:40] ^ 9);
  assign w165[68] = |(datain[39:36] ^ 14);
  assign w165[69] = |(datain[35:32] ^ 8);
  assign w165[70] = |(datain[31:28] ^ 0);
  assign w165[71] = |(datain[27:24] ^ 6);
  assign w165[72] = |(datain[23:20] ^ 0);
  assign w165[73] = |(datain[19:16] ^ 0);
  assign w165[74] = |(datain[15:12] ^ 11);
  assign w165[75] = |(datain[11:8] ^ 4);
  assign comp[165] = ~(|w165);
  wire [30-1:0] w166;
  assign w166[0] = |(datain[311:308] ^ 15);
  assign w166[1] = |(datain[307:304] ^ 15);
  assign w166[2] = |(datain[303:300] ^ 12);
  assign w166[3] = |(datain[299:296] ^ 13);
  assign w166[4] = |(datain[295:292] ^ 2);
  assign w166[5] = |(datain[291:288] ^ 1);
  assign w166[6] = |(datain[287:284] ^ 3);
  assign w166[7] = |(datain[283:280] ^ 13);
  assign w166[8] = |(datain[279:276] ^ 0);
  assign w166[9] = |(datain[275:272] ^ 1);
  assign w166[10] = |(datain[271:268] ^ 0);
  assign w166[11] = |(datain[267:264] ^ 1);
  assign w166[12] = |(datain[263:260] ^ 7);
  assign w166[13] = |(datain[259:256] ^ 4);
  assign w166[14] = |(datain[255:252] ^ 3);
  assign w166[15] = |(datain[251:248] ^ 11);
  assign w166[16] = |(datain[247:244] ^ 0);
  assign w166[17] = |(datain[243:240] ^ 6);
  assign w166[18] = |(datain[239:236] ^ 11);
  assign w166[19] = |(datain[235:232] ^ 8);
  assign w166[20] = |(datain[231:228] ^ 15);
  assign w166[21] = |(datain[227:224] ^ 1);
  assign w166[22] = |(datain[223:220] ^ 3);
  assign w166[23] = |(datain[219:216] ^ 5);
  assign w166[24] = |(datain[215:212] ^ 12);
  assign w166[25] = |(datain[211:208] ^ 13);
  assign w166[26] = |(datain[207:204] ^ 2);
  assign w166[27] = |(datain[203:200] ^ 1);
  assign w166[28] = |(datain[199:196] ^ 8);
  assign w166[29] = |(datain[195:192] ^ 12);
  assign comp[166] = ~(|w166);
  wire [32-1:0] w167;
  assign w167[0] = |(datain[311:308] ^ 5);
  assign w167[1] = |(datain[307:304] ^ 11);
  assign w167[2] = |(datain[303:300] ^ 8);
  assign w167[3] = |(datain[299:296] ^ 1);
  assign w167[4] = |(datain[295:292] ^ 12);
  assign w167[5] = |(datain[291:288] ^ 3);
  assign w167[6] = |(datain[287:284] ^ 1);
  assign w167[7] = |(datain[283:280] ^ 0);
  assign w167[8] = |(datain[279:276] ^ 0);
  assign w167[9] = |(datain[275:272] ^ 0);
  assign w167[10] = |(datain[271:268] ^ 11);
  assign w167[11] = |(datain[267:264] ^ 9);
  assign w167[12] = |(datain[263:260] ^ 9);
  assign w167[13] = |(datain[259:256] ^ 15);
  assign w167[14] = |(datain[255:252] ^ 0);
  assign w167[15] = |(datain[251:248] ^ 6);
  assign w167[16] = |(datain[247:244] ^ 3);
  assign w167[17] = |(datain[243:240] ^ 3);
  assign w167[18] = |(datain[239:236] ^ 15);
  assign w167[19] = |(datain[235:232] ^ 6);
  assign w167[20] = |(datain[231:228] ^ 8);
  assign w167[21] = |(datain[227:224] ^ 0);
  assign w167[22] = |(datain[223:220] ^ 3);
  assign w167[23] = |(datain[219:216] ^ 0);
  assign w167[24] = |(datain[215:212] ^ 5);
  assign w167[25] = |(datain[211:208] ^ 12);
  assign w167[26] = |(datain[207:204] ^ 4);
  assign w167[27] = |(datain[203:200] ^ 6);
  assign w167[28] = |(datain[199:196] ^ 14);
  assign w167[29] = |(datain[195:192] ^ 2);
  assign w167[30] = |(datain[191:188] ^ 15);
  assign w167[31] = |(datain[187:184] ^ 10);
  assign comp[167] = ~(|w167);
  wire [74-1:0] w168;
  assign w168[0] = |(datain[311:308] ^ 3);
  assign w168[1] = |(datain[307:304] ^ 3);
  assign w168[2] = |(datain[303:300] ^ 12);
  assign w168[3] = |(datain[299:296] ^ 9);
  assign w168[4] = |(datain[295:292] ^ 11);
  assign w168[5] = |(datain[291:288] ^ 8);
  assign w168[6] = |(datain[287:284] ^ 0);
  assign w168[7] = |(datain[283:280] ^ 0);
  assign w168[8] = |(datain[279:276] ^ 4);
  assign w168[9] = |(datain[275:272] ^ 2);
  assign w168[10] = |(datain[271:268] ^ 12);
  assign w168[11] = |(datain[267:264] ^ 13);
  assign w168[12] = |(datain[263:260] ^ 2);
  assign w168[13] = |(datain[259:256] ^ 1);
  assign w168[14] = |(datain[255:252] ^ 11);
  assign w168[15] = |(datain[251:248] ^ 9);
  assign w168[16] = |(datain[247:244] ^ 1);
  assign w168[17] = |(datain[243:240] ^ 12);
  assign w168[18] = |(datain[239:236] ^ 0);
  assign w168[19] = |(datain[235:232] ^ 0);
  assign w168[20] = |(datain[231:228] ^ 11);
  assign w168[21] = |(datain[227:224] ^ 10);
  assign w168[22] = |(datain[223:220] ^ 10);
  assign w168[23] = |(datain[219:216] ^ 1);
  assign w168[24] = |(datain[215:212] ^ 0);
  assign w168[25] = |(datain[211:208] ^ 2);
  assign w168[26] = |(datain[207:204] ^ 11);
  assign w168[27] = |(datain[203:200] ^ 4);
  assign w168[28] = |(datain[199:196] ^ 4);
  assign w168[29] = |(datain[195:192] ^ 0);
  assign w168[30] = |(datain[191:188] ^ 12);
  assign w168[31] = |(datain[187:184] ^ 13);
  assign w168[32] = |(datain[183:180] ^ 2);
  assign w168[33] = |(datain[179:176] ^ 1);
  assign w168[34] = |(datain[175:172] ^ 14);
  assign w168[35] = |(datain[171:168] ^ 9);
  assign w168[36] = |(datain[167:164] ^ 2);
  assign w168[37] = |(datain[163:160] ^ 4);
  assign w168[38] = |(datain[159:156] ^ 15);
  assign w168[39] = |(datain[155:152] ^ 15);
  assign w168[40] = |(datain[151:148] ^ 5);
  assign w168[41] = |(datain[147:144] ^ 11);
  assign w168[42] = |(datain[143:140] ^ 4);
  assign w168[43] = |(datain[139:136] ^ 2);
  assign w168[44] = |(datain[135:132] ^ 4);
  assign w168[45] = |(datain[131:128] ^ 5);
  assign w168[46] = |(datain[127:124] ^ 4);
  assign w168[47] = |(datain[123:120] ^ 1);
  assign w168[48] = |(datain[119:116] ^ 5);
  assign w168[49] = |(datain[115:112] ^ 6);
  assign w168[50] = |(datain[111:108] ^ 4);
  assign w168[51] = |(datain[107:104] ^ 9);
  assign w168[52] = |(datain[103:100] ^ 5);
  assign w168[53] = |(datain[99:96] ^ 3);
  assign w168[54] = |(datain[95:92] ^ 5);
  assign w168[55] = |(datain[91:88] ^ 13);
  assign w168[56] = |(datain[87:84] ^ 2);
  assign w168[57] = |(datain[83:80] ^ 0);
  assign w168[58] = |(datain[79:76] ^ 6);
  assign w168[59] = |(datain[75:72] ^ 2);
  assign w168[60] = |(datain[71:68] ^ 7);
  assign w168[61] = |(datain[67:64] ^ 9);
  assign w168[62] = |(datain[63:60] ^ 2);
  assign w168[63] = |(datain[59:56] ^ 0);
  assign w168[64] = |(datain[55:52] ^ 4);
  assign w168[65] = |(datain[51:48] ^ 3);
  assign w168[66] = |(datain[47:44] ^ 7);
  assign w168[67] = |(datain[43:40] ^ 2);
  assign w168[68] = |(datain[39:36] ^ 7);
  assign w168[69] = |(datain[35:32] ^ 9);
  assign w168[70] = |(datain[31:28] ^ 7);
  assign w168[71] = |(datain[27:24] ^ 0);
  assign w168[72] = |(datain[23:20] ^ 7);
  assign w168[73] = |(datain[19:16] ^ 4);
  assign comp[168] = ~(|w168);
  wire [74-1:0] w169;
  assign w169[0] = |(datain[311:308] ^ 9);
  assign w169[1] = |(datain[307:304] ^ 15);
  assign w169[2] = |(datain[303:300] ^ 0);
  assign w169[3] = |(datain[299:296] ^ 2);
  assign w169[4] = |(datain[295:292] ^ 8);
  assign w169[5] = |(datain[291:288] ^ 3);
  assign w169[6] = |(datain[287:284] ^ 0);
  assign w169[7] = |(datain[283:280] ^ 6);
  assign w169[8] = |(datain[279:276] ^ 9);
  assign w169[9] = |(datain[275:272] ^ 11);
  assign w169[10] = |(datain[271:268] ^ 0);
  assign w169[11] = |(datain[267:264] ^ 2);
  assign w169[12] = |(datain[263:260] ^ 2);
  assign w169[13] = |(datain[259:256] ^ 12);
  assign w169[14] = |(datain[255:252] ^ 9);
  assign w169[15] = |(datain[251:248] ^ 0);
  assign w169[16] = |(datain[247:244] ^ 11);
  assign w169[17] = |(datain[243:240] ^ 9);
  assign w169[18] = |(datain[239:236] ^ 9);
  assign w169[19] = |(datain[235:232] ^ 1);
  assign w169[20] = |(datain[231:228] ^ 0);
  assign w169[21] = |(datain[227:224] ^ 2);
  assign w169[22] = |(datain[223:220] ^ 3);
  assign w169[23] = |(datain[219:216] ^ 3);
  assign w169[24] = |(datain[215:212] ^ 13);
  assign w169[25] = |(datain[211:208] ^ 2);
  assign w169[26] = |(datain[207:204] ^ 11);
  assign w169[27] = |(datain[203:200] ^ 4);
  assign w169[28] = |(datain[199:196] ^ 4);
  assign w169[29] = |(datain[195:192] ^ 0);
  assign w169[30] = |(datain[191:188] ^ 12);
  assign w169[31] = |(datain[187:184] ^ 13);
  assign w169[32] = |(datain[183:180] ^ 2);
  assign w169[33] = |(datain[179:176] ^ 1);
  assign w169[34] = |(datain[175:172] ^ 14);
  assign w169[35] = |(datain[171:168] ^ 8);
  assign w169[36] = |(datain[167:164] ^ 2);
  assign w169[37] = |(datain[163:160] ^ 3);
  assign w169[38] = |(datain[159:156] ^ 15);
  assign w169[39] = |(datain[155:152] ^ 14);
  assign w169[40] = |(datain[151:148] ^ 11);
  assign w169[41] = |(datain[147:144] ^ 9);
  assign w169[42] = |(datain[143:140] ^ 0);
  assign w169[43] = |(datain[139:136] ^ 0);
  assign w169[44] = |(datain[135:132] ^ 0);
  assign w169[45] = |(datain[131:128] ^ 2);
  assign w169[46] = |(datain[127:124] ^ 15);
  assign w169[47] = |(datain[123:120] ^ 7);
  assign w169[48] = |(datain[119:116] ^ 15);
  assign w169[49] = |(datain[115:112] ^ 1);
  assign w169[50] = |(datain[111:108] ^ 8);
  assign w169[51] = |(datain[107:104] ^ 3);
  assign w169[52] = |(datain[103:100] ^ 15);
  assign w169[53] = |(datain[99:96] ^ 10);
  assign w169[54] = |(datain[95:92] ^ 0);
  assign w169[55] = |(datain[91:88] ^ 0);
  assign w169[56] = |(datain[87:84] ^ 7);
  assign w169[57] = |(datain[83:80] ^ 4);
  assign w169[58] = |(datain[79:76] ^ 0);
  assign w169[59] = |(datain[75:72] ^ 1);
  assign w169[60] = |(datain[71:68] ^ 4);
  assign w169[61] = |(datain[67:64] ^ 0);
  assign w169[62] = |(datain[63:60] ^ 10);
  assign w169[63] = |(datain[59:56] ^ 3);
  assign w169[64] = |(datain[55:52] ^ 9);
  assign w169[65] = |(datain[51:48] ^ 5);
  assign w169[66] = |(datain[47:44] ^ 0);
  assign w169[67] = |(datain[43:40] ^ 2);
  assign w169[68] = |(datain[39:36] ^ 8);
  assign w169[69] = |(datain[35:32] ^ 9);
  assign w169[70] = |(datain[31:28] ^ 1);
  assign w169[71] = |(datain[27:24] ^ 6);
  assign w169[72] = |(datain[23:20] ^ 9);
  assign w169[73] = |(datain[19:16] ^ 3);
  assign comp[169] = ~(|w169);
  wire [32-1:0] w170;
  assign w170[0] = |(datain[311:308] ^ 8);
  assign w170[1] = |(datain[307:304] ^ 6);
  assign w170[2] = |(datain[303:300] ^ 0);
  assign w170[3] = |(datain[299:296] ^ 0);
  assign w170[4] = |(datain[295:292] ^ 8);
  assign w170[5] = |(datain[291:288] ^ 14);
  assign w170[6] = |(datain[287:284] ^ 13);
  assign w170[7] = |(datain[283:280] ^ 11);
  assign w170[8] = |(datain[279:276] ^ 12);
  assign w170[9] = |(datain[275:272] ^ 6);
  assign w170[10] = |(datain[271:268] ^ 0);
  assign w170[11] = |(datain[267:264] ^ 6);
  assign w170[12] = |(datain[263:260] ^ 5);
  assign w170[13] = |(datain[259:256] ^ 0);
  assign w170[14] = |(datain[255:252] ^ 0);
  assign w170[15] = |(datain[251:248] ^ 7);
  assign w170[16] = |(datain[247:244] ^ 0);
  assign w170[17] = |(datain[243:240] ^ 0);
  assign w170[18] = |(datain[239:236] ^ 12);
  assign w170[19] = |(datain[235:232] ^ 6);
  assign w170[20] = |(datain[231:228] ^ 0);
  assign w170[21] = |(datain[227:224] ^ 6);
  assign w170[22] = |(datain[223:220] ^ 5);
  assign w170[23] = |(datain[219:216] ^ 1);
  assign w170[24] = |(datain[215:212] ^ 0);
  assign w170[25] = |(datain[211:208] ^ 7);
  assign w170[26] = |(datain[207:204] ^ 0);
  assign w170[27] = |(datain[203:200] ^ 0);
  assign w170[28] = |(datain[199:196] ^ 10);
  assign w170[29] = |(datain[195:192] ^ 3);
  assign w170[30] = |(datain[191:188] ^ 3);
  assign w170[31] = |(datain[187:184] ^ 11);
  assign comp[170] = ~(|w170);
  wire [30-1:0] w171;
  assign w171[0] = |(datain[311:308] ^ 12);
  assign w171[1] = |(datain[307:304] ^ 0);
  assign w171[2] = |(datain[303:300] ^ 3);
  assign w171[3] = |(datain[299:296] ^ 3);
  assign w171[4] = |(datain[295:292] ^ 15);
  assign w171[5] = |(datain[291:288] ^ 15);
  assign w171[6] = |(datain[287:284] ^ 3);
  assign w171[7] = |(datain[283:280] ^ 3);
  assign w171[8] = |(datain[279:276] ^ 12);
  assign w171[9] = |(datain[275:272] ^ 0);
  assign w171[10] = |(datain[271:268] ^ 11);
  assign w171[11] = |(datain[267:264] ^ 9);
  assign w171[12] = |(datain[263:260] ^ 15);
  assign w171[13] = |(datain[259:256] ^ 15);
  assign w171[14] = |(datain[255:252] ^ 7);
  assign w171[15] = |(datain[251:248] ^ 15);
  assign w171[16] = |(datain[247:244] ^ 15);
  assign w171[17] = |(datain[243:240] ^ 12);
  assign w171[18] = |(datain[239:236] ^ 15);
  assign w171[19] = |(datain[235:232] ^ 2);
  assign w171[20] = |(datain[231:228] ^ 10);
  assign w171[21] = |(datain[227:224] ^ 14);
  assign w171[22] = |(datain[223:220] ^ 2);
  assign w171[23] = |(datain[219:216] ^ 6);
  assign w171[24] = |(datain[215:212] ^ 15);
  assign w171[25] = |(datain[211:208] ^ 6);
  assign w171[26] = |(datain[207:204] ^ 0);
  assign w171[27] = |(datain[203:200] ^ 5);
  assign w171[28] = |(datain[199:196] ^ 15);
  assign w171[29] = |(datain[195:192] ^ 15);
  assign comp[171] = ~(|w171);
  wire [38-1:0] w172;
  assign w172[0] = |(datain[311:308] ^ 0);
  assign w172[1] = |(datain[307:304] ^ 2);
  assign w172[2] = |(datain[303:300] ^ 0);
  assign w172[3] = |(datain[299:296] ^ 0);
  assign w172[4] = |(datain[295:292] ^ 11);
  assign w172[5] = |(datain[291:288] ^ 4);
  assign w172[6] = |(datain[287:284] ^ 3);
  assign w172[7] = |(datain[283:280] ^ 15);
  assign w172[8] = |(datain[279:276] ^ 12);
  assign w172[9] = |(datain[275:272] ^ 13);
  assign w172[10] = |(datain[271:268] ^ 2);
  assign w172[11] = |(datain[267:264] ^ 1);
  assign w172[12] = |(datain[263:260] ^ 8);
  assign w172[13] = |(datain[259:256] ^ 1);
  assign w172[14] = |(datain[255:252] ^ 3);
  assign w172[15] = |(datain[251:248] ^ 13);
  assign w172[16] = |(datain[247:244] ^ 0);
  assign w172[17] = |(datain[243:240] ^ 7);
  assign w172[18] = |(datain[239:236] ^ 0);
  assign w172[19] = |(datain[235:232] ^ 8);
  assign w172[20] = |(datain[231:228] ^ 7);
  assign w172[21] = |(datain[227:224] ^ 4);
  assign w172[22] = |(datain[223:220] ^ 13);
  assign w172[23] = |(datain[219:216] ^ 15);
  assign w172[24] = |(datain[215:212] ^ 3);
  assign w172[25] = |(datain[211:208] ^ 3);
  assign w172[26] = |(datain[207:204] ^ 12);
  assign w172[27] = |(datain[203:200] ^ 9);
  assign w172[28] = |(datain[199:196] ^ 11);
  assign w172[29] = |(datain[195:192] ^ 8);
  assign w172[30] = |(datain[191:188] ^ 0);
  assign w172[31] = |(datain[187:184] ^ 2);
  assign w172[32] = |(datain[183:180] ^ 4);
  assign w172[33] = |(datain[179:176] ^ 2);
  assign w172[34] = |(datain[175:172] ^ 12);
  assign w172[35] = |(datain[171:168] ^ 13);
  assign w172[36] = |(datain[167:164] ^ 2);
  assign w172[37] = |(datain[163:160] ^ 1);
  assign comp[172] = ~(|w172);
  wire [32-1:0] w173;
  assign w173[0] = |(datain[311:308] ^ 8);
  assign w173[1] = |(datain[307:304] ^ 11);
  assign w173[2] = |(datain[303:300] ^ 13);
  assign w173[3] = |(datain[299:296] ^ 7);
  assign w173[4] = |(datain[295:292] ^ 11);
  assign w173[5] = |(datain[291:288] ^ 9);
  assign w173[6] = |(datain[287:284] ^ 0);
  assign w173[7] = |(datain[283:280] ^ 2);
  assign w173[8] = |(datain[279:276] ^ 0);
  assign w173[9] = |(datain[275:272] ^ 0);
  assign w173[10] = |(datain[271:268] ^ 11);
  assign w173[11] = |(datain[267:264] ^ 4);
  assign w173[12] = |(datain[263:260] ^ 3);
  assign w173[13] = |(datain[259:256] ^ 15);
  assign w173[14] = |(datain[255:252] ^ 12);
  assign w173[15] = |(datain[251:248] ^ 13);
  assign w173[16] = |(datain[247:244] ^ 2);
  assign w173[17] = |(datain[243:240] ^ 1);
  assign w173[18] = |(datain[239:236] ^ 8);
  assign w173[19] = |(datain[235:232] ^ 1);
  assign w173[20] = |(datain[231:228] ^ 3);
  assign w173[21] = |(datain[227:224] ^ 13);
  assign w173[22] = |(datain[223:220] ^ 0);
  assign w173[23] = |(datain[219:216] ^ 7);
  assign w173[24] = |(datain[215:212] ^ 0);
  assign w173[25] = |(datain[211:208] ^ 8);
  assign w173[26] = |(datain[207:204] ^ 7);
  assign w173[27] = |(datain[203:200] ^ 4);
  assign w173[28] = |(datain[199:196] ^ 13);
  assign w173[29] = |(datain[195:192] ^ 15);
  assign w173[30] = |(datain[191:188] ^ 3);
  assign w173[31] = |(datain[187:184] ^ 3);
  assign comp[173] = ~(|w173);
  wire [28-1:0] w174;
  assign w174[0] = |(datain[311:308] ^ 0);
  assign w174[1] = |(datain[307:304] ^ 5);
  assign w174[2] = |(datain[303:300] ^ 0);
  assign w174[3] = |(datain[299:296] ^ 0);
  assign w174[4] = |(datain[295:292] ^ 12);
  assign w174[5] = |(datain[291:288] ^ 13);
  assign w174[6] = |(datain[287:284] ^ 2);
  assign w174[7] = |(datain[283:280] ^ 15);
  assign w174[8] = |(datain[279:276] ^ 5);
  assign w174[9] = |(datain[275:272] ^ 3);
  assign w174[10] = |(datain[271:268] ^ 4);
  assign w174[11] = |(datain[267:264] ^ 11);
  assign w174[12] = |(datain[263:260] ^ 4);
  assign w174[13] = |(datain[259:256] ^ 11);
  assign w174[14] = |(datain[255:252] ^ 2);
  assign w174[15] = |(datain[251:248] ^ 6);
  assign w174[16] = |(datain[247:244] ^ 8);
  assign w174[17] = |(datain[243:240] ^ 8);
  assign w174[18] = |(datain[239:236] ^ 1);
  assign w174[19] = |(datain[235:232] ^ 13);
  assign w174[20] = |(datain[231:228] ^ 11);
  assign w174[21] = |(datain[227:224] ^ 8);
  assign w174[22] = |(datain[223:220] ^ 1);
  assign w174[23] = |(datain[219:216] ^ 6);
  assign w174[24] = |(datain[215:212] ^ 1);
  assign w174[25] = |(datain[211:208] ^ 2);
  assign w174[26] = |(datain[207:204] ^ 12);
  assign w174[27] = |(datain[203:200] ^ 13);
  assign comp[174] = ~(|w174);
  wire [46-1:0] w175;
  assign w175[0] = |(datain[311:308] ^ 2);
  assign w175[1] = |(datain[307:304] ^ 0);
  assign w175[2] = |(datain[303:300] ^ 1);
  assign w175[3] = |(datain[299:296] ^ 2);
  assign w175[4] = |(datain[295:292] ^ 11);
  assign w175[5] = |(datain[291:288] ^ 11);
  assign w175[6] = |(datain[287:284] ^ 0);
  assign w175[7] = |(datain[283:280] ^ 5);
  assign w175[8] = |(datain[279:276] ^ 0);
  assign w175[9] = |(datain[275:272] ^ 0);
  assign w175[10] = |(datain[271:268] ^ 12);
  assign w175[11] = |(datain[267:264] ^ 13);
  assign w175[12] = |(datain[263:260] ^ 2);
  assign w175[13] = |(datain[259:256] ^ 15);
  assign w175[14] = |(datain[255:252] ^ 5);
  assign w175[15] = |(datain[251:248] ^ 3);
  assign w175[16] = |(datain[247:244] ^ 4);
  assign w175[17] = |(datain[243:240] ^ 11);
  assign w175[18] = |(datain[239:236] ^ 4);
  assign w175[19] = |(datain[235:232] ^ 11);
  assign w175[20] = |(datain[231:228] ^ 2);
  assign w175[21] = |(datain[227:224] ^ 6);
  assign w175[22] = |(datain[223:220] ^ 8);
  assign w175[23] = |(datain[219:216] ^ 8);
  assign w175[24] = |(datain[215:212] ^ 1);
  assign w175[25] = |(datain[211:208] ^ 13);
  assign w175[26] = |(datain[207:204] ^ 11);
  assign w175[27] = |(datain[203:200] ^ 8);
  assign w175[28] = |(datain[199:196] ^ 1);
  assign w175[29] = |(datain[195:192] ^ 6);
  assign w175[30] = |(datain[191:188] ^ 1);
  assign w175[31] = |(datain[187:184] ^ 2);
  assign w175[32] = |(datain[183:180] ^ 12);
  assign w175[33] = |(datain[179:176] ^ 13);
  assign w175[34] = |(datain[175:172] ^ 2);
  assign w175[35] = |(datain[171:168] ^ 15);
  assign w175[36] = |(datain[167:164] ^ 4);
  assign w175[37] = |(datain[163:160] ^ 11);
  assign w175[38] = |(datain[159:156] ^ 4);
  assign w175[39] = |(datain[155:152] ^ 11);
  assign w175[40] = |(datain[151:148] ^ 2);
  assign w175[41] = |(datain[147:144] ^ 6);
  assign w175[42] = |(datain[143:140] ^ 8);
  assign w175[43] = |(datain[139:136] ^ 9);
  assign w175[44] = |(datain[135:132] ^ 1);
  assign w175[45] = |(datain[131:128] ^ 13);
  assign comp[175] = ~(|w175);
  wire [32-1:0] w176;
  assign w176[0] = |(datain[311:308] ^ 1);
  assign w176[1] = |(datain[307:304] ^ 14);
  assign w176[2] = |(datain[303:300] ^ 11);
  assign w176[3] = |(datain[299:296] ^ 8);
  assign w176[4] = |(datain[295:292] ^ 0);
  assign w176[5] = |(datain[291:288] ^ 3);
  assign w176[6] = |(datain[287:284] ^ 1);
  assign w176[7] = |(datain[283:280] ^ 2);
  assign w176[8] = |(datain[279:276] ^ 12);
  assign w176[9] = |(datain[275:272] ^ 13);
  assign w176[10] = |(datain[271:268] ^ 2);
  assign w176[11] = |(datain[267:264] ^ 15);
  assign w176[12] = |(datain[263:260] ^ 2);
  assign w176[13] = |(datain[259:256] ^ 14);
  assign w176[14] = |(datain[255:252] ^ 8);
  assign w176[15] = |(datain[251:248] ^ 12);
  assign w176[16] = |(datain[247:244] ^ 1);
  assign w176[17] = |(datain[243:240] ^ 14);
  assign w176[18] = |(datain[239:236] ^ 0);
  assign w176[19] = |(datain[235:232] ^ 4);
  assign w176[20] = |(datain[231:228] ^ 0);
  assign w176[21] = |(datain[227:224] ^ 9);
  assign w176[22] = |(datain[223:220] ^ 3);
  assign w176[23] = |(datain[219:216] ^ 3);
  assign w176[24] = |(datain[215:212] ^ 15);
  assign w176[25] = |(datain[211:208] ^ 6);
  assign w176[26] = |(datain[207:204] ^ 8);
  assign w176[27] = |(datain[203:200] ^ 14);
  assign w176[28] = |(datain[199:196] ^ 13);
  assign w176[29] = |(datain[195:192] ^ 14);
  assign w176[30] = |(datain[191:188] ^ 11);
  assign w176[31] = |(datain[187:184] ^ 15);
  assign comp[176] = ~(|w176);
  wire [46-1:0] w177;
  assign w177[0] = |(datain[311:308] ^ 12);
  assign w177[1] = |(datain[307:304] ^ 0);
  assign w177[2] = |(datain[303:300] ^ 3);
  assign w177[3] = |(datain[299:296] ^ 3);
  assign w177[4] = |(datain[295:292] ^ 15);
  assign w177[5] = |(datain[291:288] ^ 15);
  assign w177[6] = |(datain[287:284] ^ 3);
  assign w177[7] = |(datain[283:280] ^ 3);
  assign w177[8] = |(datain[279:276] ^ 12);
  assign w177[9] = |(datain[275:272] ^ 0);
  assign w177[10] = |(datain[271:268] ^ 11);
  assign w177[11] = |(datain[267:264] ^ 9);
  assign w177[12] = |(datain[263:260] ^ 15);
  assign w177[13] = |(datain[259:256] ^ 15);
  assign w177[14] = |(datain[255:252] ^ 7);
  assign w177[15] = |(datain[251:248] ^ 15);
  assign w177[16] = |(datain[247:244] ^ 15);
  assign w177[17] = |(datain[243:240] ^ 12);
  assign w177[18] = |(datain[239:236] ^ 15);
  assign w177[19] = |(datain[235:232] ^ 2);
  assign w177[20] = |(datain[231:228] ^ 10);
  assign w177[21] = |(datain[227:224] ^ 14);
  assign w177[22] = |(datain[223:220] ^ 2);
  assign w177[23] = |(datain[219:216] ^ 6);
  assign w177[24] = |(datain[215:212] ^ 15);
  assign w177[25] = |(datain[211:208] ^ 6);
  assign w177[26] = |(datain[207:204] ^ 0);
  assign w177[27] = |(datain[203:200] ^ 5);
  assign w177[28] = |(datain[199:196] ^ 15);
  assign w177[29] = |(datain[195:192] ^ 15);
  assign w177[30] = |(datain[191:188] ^ 7);
  assign w177[31] = |(datain[187:184] ^ 5);
  assign w177[32] = |(datain[183:180] ^ 15);
  assign w177[33] = |(datain[179:176] ^ 8);
  assign w177[34] = |(datain[175:172] ^ 8);
  assign w177[35] = |(datain[171:168] ^ 3);
  assign w177[36] = |(datain[167:164] ^ 12);
  assign w177[37] = |(datain[163:160] ^ 7);
  assign w177[38] = |(datain[159:156] ^ 0);
  assign w177[39] = |(datain[155:152] ^ 3);
  assign w177[40] = |(datain[151:148] ^ 8);
  assign w177[41] = |(datain[147:144] ^ 11);
  assign w177[42] = |(datain[143:140] ^ 13);
  assign w177[43] = |(datain[139:136] ^ 7);
  assign w177[44] = |(datain[135:132] ^ 2);
  assign w177[45] = |(datain[131:128] ^ 14);
  assign comp[177] = ~(|w177);
  wire [28-1:0] w178;
  assign w178[0] = |(datain[311:308] ^ 0);
  assign w178[1] = |(datain[307:304] ^ 1);
  assign w178[2] = |(datain[303:300] ^ 8);
  assign w178[3] = |(datain[299:296] ^ 10);
  assign w178[4] = |(datain[295:292] ^ 2);
  assign w178[5] = |(datain[291:288] ^ 15);
  assign w178[6] = |(datain[287:284] ^ 3);
  assign w178[7] = |(datain[283:280] ^ 2);
  assign w178[8] = |(datain[279:276] ^ 2);
  assign w178[9] = |(datain[275:272] ^ 14);
  assign w178[10] = |(datain[271:268] ^ 0);
  assign w178[11] = |(datain[267:264] ^ 3);
  assign w178[12] = |(datain[263:260] ^ 0);
  assign w178[13] = |(datain[259:256] ^ 1);
  assign w178[14] = |(datain[255:252] ^ 8);
  assign w178[15] = |(datain[251:248] ^ 8);
  assign w178[16] = |(datain[247:244] ^ 2);
  assign w178[17] = |(datain[243:240] ^ 15);
  assign w178[18] = |(datain[239:236] ^ 4);
  assign w178[19] = |(datain[235:232] ^ 3);
  assign w178[20] = |(datain[231:228] ^ 8);
  assign w178[21] = |(datain[227:224] ^ 1);
  assign w178[22] = |(datain[223:220] ^ 15);
  assign w178[23] = |(datain[219:216] ^ 11);
  assign w178[24] = |(datain[215:212] ^ 0);
  assign w178[25] = |(datain[211:208] ^ 0);
  assign w178[26] = |(datain[207:204] ^ 0);
  assign w178[27] = |(datain[203:200] ^ 9);
  assign comp[178] = ~(|w178);
  wire [30-1:0] w179;
  assign w179[0] = |(datain[311:308] ^ 13);
  assign w179[1] = |(datain[307:304] ^ 2);
  assign w179[2] = |(datain[303:300] ^ 11);
  assign w179[3] = |(datain[299:296] ^ 8);
  assign w179[4] = |(datain[295:292] ^ 0);
  assign w179[5] = |(datain[291:288] ^ 0);
  assign w179[6] = |(datain[287:284] ^ 4);
  assign w179[7] = |(datain[283:280] ^ 2);
  assign w179[8] = |(datain[279:276] ^ 12);
  assign w179[9] = |(datain[275:272] ^ 13);
  assign w179[10] = |(datain[271:268] ^ 2);
  assign w179[11] = |(datain[267:264] ^ 1);
  assign w179[12] = |(datain[263:260] ^ 8);
  assign w179[13] = |(datain[259:256] ^ 11);
  assign w179[14] = |(datain[255:252] ^ 12);
  assign w179[15] = |(datain[251:248] ^ 14);
  assign w179[16] = |(datain[247:244] ^ 11);
  assign w179[17] = |(datain[243:240] ^ 4);
  assign w179[18] = |(datain[239:236] ^ 4);
  assign w179[19] = |(datain[235:232] ^ 0);
  assign w179[20] = |(datain[231:228] ^ 12);
  assign w179[21] = |(datain[227:224] ^ 13);
  assign w179[22] = |(datain[223:220] ^ 2);
  assign w179[23] = |(datain[219:216] ^ 1);
  assign w179[24] = |(datain[215:212] ^ 2);
  assign w179[25] = |(datain[211:208] ^ 14);
  assign w179[26] = |(datain[207:204] ^ 8);
  assign w179[27] = |(datain[203:200] ^ 11);
  assign w179[28] = |(datain[199:196] ^ 0);
  assign w179[29] = |(datain[195:192] ^ 14);
  assign comp[179] = ~(|w179);
  wire [74-1:0] w180;
  assign w180[0] = |(datain[311:308] ^ 12);
  assign w180[1] = |(datain[307:304] ^ 7);
  assign w180[2] = |(datain[303:300] ^ 0);
  assign w180[3] = |(datain[299:296] ^ 3);
  assign w180[4] = |(datain[295:292] ^ 11);
  assign w180[5] = |(datain[291:288] ^ 0);
  assign w180[6] = |(datain[287:284] ^ 0);
  assign w180[7] = |(datain[283:280] ^ 0);
  assign w180[8] = |(datain[279:276] ^ 14);
  assign w180[9] = |(datain[275:272] ^ 8);
  assign w180[10] = |(datain[271:268] ^ 3);
  assign w180[11] = |(datain[267:264] ^ 14);
  assign w180[12] = |(datain[263:260] ^ 15);
  assign w180[13] = |(datain[259:256] ^ 15);
  assign w180[14] = |(datain[255:252] ^ 11);
  assign w180[15] = |(datain[251:248] ^ 4);
  assign w180[16] = |(datain[247:244] ^ 4);
  assign w180[17] = |(datain[243:240] ^ 0);
  assign w180[18] = |(datain[239:236] ^ 11);
  assign w180[19] = |(datain[235:232] ^ 10);
  assign w180[20] = |(datain[231:228] ^ 14);
  assign w180[21] = |(datain[227:224] ^ 15);
  assign w180[22] = |(datain[223:220] ^ 0);
  assign w180[23] = |(datain[219:216] ^ 3);
  assign w180[24] = |(datain[215:212] ^ 11);
  assign w180[25] = |(datain[211:208] ^ 9);
  assign w180[26] = |(datain[207:204] ^ 1);
  assign w180[27] = |(datain[203:200] ^ 10);
  assign w180[28] = |(datain[199:196] ^ 0);
  assign w180[29] = |(datain[195:192] ^ 0);
  assign w180[30] = |(datain[191:188] ^ 12);
  assign w180[31] = |(datain[187:184] ^ 13);
  assign w180[32] = |(datain[183:180] ^ 2);
  assign w180[33] = |(datain[179:176] ^ 1);
  assign w180[34] = |(datain[175:172] ^ 14);
  assign w180[35] = |(datain[171:168] ^ 8);
  assign w180[36] = |(datain[167:164] ^ 2);
  assign w180[37] = |(datain[163:160] ^ 15);
  assign w180[38] = |(datain[159:156] ^ 15);
  assign w180[39] = |(datain[155:152] ^ 15);
  assign w180[40] = |(datain[151:148] ^ 8);
  assign w180[41] = |(datain[147:144] ^ 10);
  assign w180[42] = |(datain[143:140] ^ 1);
  assign w180[43] = |(datain[139:136] ^ 6);
  assign w180[44] = |(datain[135:132] ^ 0);
  assign w180[45] = |(datain[131:128] ^ 8);
  assign w180[46] = |(datain[127:124] ^ 0);
  assign w180[47] = |(datain[123:120] ^ 0);
  assign w180[48] = |(datain[119:116] ^ 10);
  assign w180[49] = |(datain[115:112] ^ 1);
  assign w180[50] = |(datain[111:108] ^ 15);
  assign w180[51] = |(datain[107:104] ^ 3);
  assign w180[52] = |(datain[103:100] ^ 0);
  assign w180[53] = |(datain[99:96] ^ 1);
  assign w180[54] = |(datain[95:92] ^ 8);
  assign w180[55] = |(datain[91:88] ^ 6);
  assign w180[56] = |(datain[87:84] ^ 2);
  assign w180[57] = |(datain[83:80] ^ 6);
  assign w180[58] = |(datain[79:76] ^ 0);
  assign w180[59] = |(datain[75:72] ^ 13);
  assign w180[60] = |(datain[71:68] ^ 0);
  assign w180[61] = |(datain[67:64] ^ 0);
  assign w180[62] = |(datain[63:60] ^ 8);
  assign w180[63] = |(datain[59:56] ^ 6);
  assign w180[64] = |(datain[55:52] ^ 14);
  assign w180[65] = |(datain[51:48] ^ 0);
  assign w180[66] = |(datain[47:44] ^ 10);
  assign w180[67] = |(datain[43:40] ^ 3);
  assign w180[68] = |(datain[39:36] ^ 15);
  assign w180[69] = |(datain[35:32] ^ 3);
  assign w180[70] = |(datain[31:28] ^ 0);
  assign w180[71] = |(datain[27:24] ^ 1);
  assign w180[72] = |(datain[23:20] ^ 10);
  assign w180[73] = |(datain[19:16] ^ 1);
  assign comp[180] = ~(|w180);
  wire [76-1:0] w181;
  assign w181[0] = |(datain[311:308] ^ 3);
  assign w181[1] = |(datain[307:304] ^ 3);
  assign w181[2] = |(datain[303:300] ^ 12);
  assign w181[3] = |(datain[299:296] ^ 9);
  assign w181[4] = |(datain[295:292] ^ 11);
  assign w181[5] = |(datain[291:288] ^ 8);
  assign w181[6] = |(datain[287:284] ^ 0);
  assign w181[7] = |(datain[283:280] ^ 0);
  assign w181[8] = |(datain[279:276] ^ 4);
  assign w181[9] = |(datain[275:272] ^ 2);
  assign w181[10] = |(datain[271:268] ^ 9);
  assign w181[11] = |(datain[267:264] ^ 9);
  assign w181[12] = |(datain[263:260] ^ 12);
  assign w181[13] = |(datain[259:256] ^ 13);
  assign w181[14] = |(datain[255:252] ^ 2);
  assign w181[15] = |(datain[251:248] ^ 1);
  assign w181[16] = |(datain[247:244] ^ 11);
  assign w181[17] = |(datain[243:240] ^ 9);
  assign w181[18] = |(datain[239:236] ^ 1);
  assign w181[19] = |(datain[235:232] ^ 10);
  assign w181[20] = |(datain[231:228] ^ 0);
  assign w181[21] = |(datain[227:224] ^ 0);
  assign w181[22] = |(datain[223:220] ^ 11);
  assign w181[23] = |(datain[219:216] ^ 10);
  assign w181[24] = |(datain[215:212] ^ 11);
  assign w181[25] = |(datain[211:208] ^ 10);
  assign w181[26] = |(datain[207:204] ^ 0);
  assign w181[27] = |(datain[203:200] ^ 1);
  assign w181[28] = |(datain[199:196] ^ 11);
  assign w181[29] = |(datain[195:192] ^ 4);
  assign w181[30] = |(datain[191:188] ^ 4);
  assign w181[31] = |(datain[187:184] ^ 0);
  assign w181[32] = |(datain[183:180] ^ 12);
  assign w181[33] = |(datain[179:176] ^ 13);
  assign w181[34] = |(datain[175:172] ^ 2);
  assign w181[35] = |(datain[171:168] ^ 1);
  assign w181[36] = |(datain[167:164] ^ 11);
  assign w181[37] = |(datain[163:160] ^ 8);
  assign w181[38] = |(datain[159:156] ^ 0);
  assign w181[39] = |(datain[155:152] ^ 1);
  assign w181[40] = |(datain[151:148] ^ 5);
  assign w181[41] = |(datain[147:144] ^ 7);
  assign w181[42] = |(datain[143:140] ^ 5);
  assign w181[43] = |(datain[139:136] ^ 10);
  assign w181[44] = |(datain[135:132] ^ 5);
  assign w181[45] = |(datain[131:128] ^ 9);
  assign w181[46] = |(datain[127:124] ^ 12);
  assign w181[47] = |(datain[123:120] ^ 13);
  assign w181[48] = |(datain[119:116] ^ 2);
  assign w181[49] = |(datain[115:112] ^ 1);
  assign w181[50] = |(datain[111:108] ^ 11);
  assign w181[51] = |(datain[107:104] ^ 4);
  assign w181[52] = |(datain[103:100] ^ 3);
  assign w181[53] = |(datain[99:96] ^ 14);
  assign w181[54] = |(datain[95:92] ^ 12);
  assign w181[55] = |(datain[91:88] ^ 13);
  assign w181[56] = |(datain[87:84] ^ 2);
  assign w181[57] = |(datain[83:80] ^ 1);
  assign w181[58] = |(datain[79:76] ^ 5);
  assign w181[59] = |(datain[75:72] ^ 8);
  assign w181[60] = |(datain[71:68] ^ 5);
  assign w181[61] = |(datain[67:64] ^ 10);
  assign w181[62] = |(datain[63:60] ^ 1);
  assign w181[63] = |(datain[59:56] ^ 15);
  assign w181[64] = |(datain[55:52] ^ 5);
  assign w181[65] = |(datain[51:48] ^ 9);
  assign w181[66] = |(datain[47:44] ^ 12);
  assign w181[67] = |(datain[43:40] ^ 13);
  assign w181[68] = |(datain[39:36] ^ 2);
  assign w181[69] = |(datain[35:32] ^ 1);
  assign w181[70] = |(datain[31:28] ^ 5);
  assign w181[71] = |(datain[27:24] ^ 10);
  assign w181[72] = |(datain[23:20] ^ 1);
  assign w181[73] = |(datain[19:16] ^ 15);
  assign w181[74] = |(datain[15:12] ^ 11);
  assign w181[75] = |(datain[11:8] ^ 8);
  assign comp[181] = ~(|w181);
  wire [28-1:0] w182;
  assign w182[0] = |(datain[311:308] ^ 0);
  assign w182[1] = |(datain[307:304] ^ 3);
  assign w182[2] = |(datain[303:300] ^ 0);
  assign w182[3] = |(datain[299:296] ^ 1);
  assign w182[4] = |(datain[295:292] ^ 0);
  assign w182[5] = |(datain[291:288] ^ 1);
  assign w182[6] = |(datain[287:284] ^ 12);
  assign w182[7] = |(datain[283:280] ^ 6);
  assign w182[8] = |(datain[279:276] ^ 11);
  assign w182[9] = |(datain[275:272] ^ 9);
  assign w182[10] = |(datain[271:268] ^ 0);
  assign w182[11] = |(datain[267:264] ^ 4);
  assign w182[12] = |(datain[263:260] ^ 0);
  assign w182[13] = |(datain[259:256] ^ 0);
  assign w182[14] = |(datain[255:252] ^ 8);
  assign w182[15] = |(datain[251:248] ^ 12);
  assign w182[16] = |(datain[247:244] ^ 12);
  assign w182[17] = |(datain[243:240] ^ 8);
  assign w182[18] = |(datain[239:236] ^ 8);
  assign w182[19] = |(datain[235:232] ^ 14);
  assign w182[20] = |(datain[231:228] ^ 12);
  assign w182[21] = |(datain[227:224] ^ 0);
  assign w182[22] = |(datain[223:220] ^ 8);
  assign w182[23] = |(datain[219:216] ^ 14);
  assign w182[24] = |(datain[215:212] ^ 13);
  assign w182[25] = |(datain[211:208] ^ 8);
  assign w182[26] = |(datain[207:204] ^ 8);
  assign w182[27] = |(datain[203:200] ^ 15);
  assign comp[182] = ~(|w182);
  wire [32-1:0] w183;
  assign w183[0] = |(datain[311:308] ^ 0);
  assign w183[1] = |(datain[307:304] ^ 1);
  assign w183[2] = |(datain[303:300] ^ 8);
  assign w183[3] = |(datain[299:296] ^ 9);
  assign w183[4] = |(datain[295:292] ^ 0);
  assign w183[5] = |(datain[291:288] ^ 4);
  assign w183[6] = |(datain[287:284] ^ 11);
  assign w183[7] = |(datain[283:280] ^ 4);
  assign w183[8] = |(datain[279:276] ^ 4);
  assign w183[9] = |(datain[275:272] ^ 0);
  assign w183[10] = |(datain[271:268] ^ 8);
  assign w183[11] = |(datain[267:264] ^ 11);
  assign w183[12] = |(datain[263:260] ^ 13);
  assign w183[13] = |(datain[259:256] ^ 7);
  assign w183[14] = |(datain[255:252] ^ 8);
  assign w183[15] = |(datain[251:248] ^ 1);
  assign w183[16] = |(datain[247:244] ^ 12);
  assign w183[17] = |(datain[243:240] ^ 2);
  assign w183[18] = |(datain[239:236] ^ 0);
  assign w183[19] = |(datain[235:232] ^ 3);
  assign w183[20] = |(datain[231:228] ^ 0);
  assign w183[21] = |(datain[227:224] ^ 1);
  assign w183[22] = |(datain[223:220] ^ 11);
  assign w183[23] = |(datain[219:216] ^ 9);
  assign w183[24] = |(datain[215:212] ^ 11);
  assign w183[25] = |(datain[211:208] ^ 0);
  assign w183[26] = |(datain[207:204] ^ 0);
  assign w183[27] = |(datain[203:200] ^ 9);
  assign w183[28] = |(datain[199:196] ^ 12);
  assign w183[29] = |(datain[195:192] ^ 13);
  assign w183[30] = |(datain[191:188] ^ 2);
  assign w183[31] = |(datain[187:184] ^ 1);
  assign comp[183] = ~(|w183);
  wire [30-1:0] w184;
  assign w184[0] = |(datain[311:308] ^ 5);
  assign w184[1] = |(datain[307:304] ^ 14);
  assign w184[2] = |(datain[303:300] ^ 14);
  assign w184[3] = |(datain[299:296] ^ 9);
  assign w184[4] = |(datain[295:292] ^ 4);
  assign w184[5] = |(datain[291:288] ^ 6);
  assign w184[6] = |(datain[287:284] ^ 0);
  assign w184[7] = |(datain[283:280] ^ 0);
  assign w184[8] = |(datain[279:276] ^ 5);
  assign w184[9] = |(datain[275:272] ^ 14);
  assign w184[10] = |(datain[271:268] ^ 11);
  assign w184[11] = |(datain[267:264] ^ 4);
  assign w184[12] = |(datain[263:260] ^ 3);
  assign w184[13] = |(datain[259:256] ^ 13);
  assign w184[14] = |(datain[255:252] ^ 11);
  assign w184[15] = |(datain[251:248] ^ 0);
  assign w184[16] = |(datain[247:244] ^ 0);
  assign w184[17] = |(datain[243:240] ^ 2);
  assign w184[18] = |(datain[239:236] ^ 8);
  assign w184[19] = |(datain[235:232] ^ 11);
  assign w184[20] = |(datain[231:228] ^ 13);
  assign w184[21] = |(datain[227:224] ^ 6);
  assign w184[22] = |(datain[223:220] ^ 8);
  assign w184[23] = |(datain[219:216] ^ 1);
  assign w184[24] = |(datain[215:212] ^ 12);
  assign w184[25] = |(datain[211:208] ^ 2);
  assign w184[26] = |(datain[207:204] ^ 1);
  assign w184[27] = |(datain[203:200] ^ 14);
  assign w184[28] = |(datain[199:196] ^ 0);
  assign w184[29] = |(datain[195:192] ^ 0);
  assign comp[184] = ~(|w184);
  wire [30-1:0] w185;
  assign w185[0] = |(datain[311:308] ^ 12);
  assign w185[1] = |(datain[307:304] ^ 6);
  assign w185[2] = |(datain[303:300] ^ 0);
  assign w185[3] = |(datain[299:296] ^ 3);
  assign w185[4] = |(datain[295:292] ^ 0);
  assign w185[5] = |(datain[291:288] ^ 1);
  assign w185[6] = |(datain[287:284] ^ 0);
  assign w185[7] = |(datain[283:280] ^ 1);
  assign w185[8] = |(datain[279:276] ^ 12);
  assign w185[9] = |(datain[275:272] ^ 6);
  assign w185[10] = |(datain[271:268] ^ 11);
  assign w185[11] = |(datain[267:264] ^ 9);
  assign w185[12] = |(datain[263:260] ^ 0);
  assign w185[13] = |(datain[259:256] ^ 4);
  assign w185[14] = |(datain[255:252] ^ 0);
  assign w185[15] = |(datain[251:248] ^ 0);
  assign w185[16] = |(datain[247:244] ^ 8);
  assign w185[17] = |(datain[243:240] ^ 12);
  assign w185[18] = |(datain[239:236] ^ 12);
  assign w185[19] = |(datain[235:232] ^ 8);
  assign w185[20] = |(datain[231:228] ^ 8);
  assign w185[21] = |(datain[227:224] ^ 14);
  assign w185[22] = |(datain[223:220] ^ 12);
  assign w185[23] = |(datain[219:216] ^ 0);
  assign w185[24] = |(datain[215:212] ^ 8);
  assign w185[25] = |(datain[211:208] ^ 14);
  assign w185[26] = |(datain[207:204] ^ 13);
  assign w185[27] = |(datain[203:200] ^ 8);
  assign w185[28] = |(datain[199:196] ^ 11);
  assign w185[29] = |(datain[195:192] ^ 15);
  assign comp[185] = ~(|w185);
  wire [32-1:0] w186;
  assign w186[0] = |(datain[311:308] ^ 11);
  assign w186[1] = |(datain[307:304] ^ 4);
  assign w186[2] = |(datain[303:300] ^ 2);
  assign w186[3] = |(datain[299:296] ^ 10);
  assign w186[4] = |(datain[295:292] ^ 12);
  assign w186[5] = |(datain[291:288] ^ 13);
  assign w186[6] = |(datain[287:284] ^ 2);
  assign w186[7] = |(datain[283:280] ^ 1);
  assign w186[8] = |(datain[279:276] ^ 8);
  assign w186[9] = |(datain[275:272] ^ 1);
  assign w186[10] = |(datain[271:268] ^ 15);
  assign w186[11] = |(datain[267:264] ^ 9);
  assign w186[12] = |(datain[263:260] ^ 12);
  assign w186[13] = |(datain[259:256] ^ 4);
  assign w186[14] = |(datain[255:252] ^ 0);
  assign w186[15] = |(datain[251:248] ^ 7);
  assign w186[16] = |(datain[247:244] ^ 7);
  assign w186[17] = |(datain[243:240] ^ 2);
  assign w186[18] = |(datain[239:236] ^ 0);
  assign w186[19] = |(datain[235:232] ^ 8);
  assign w186[20] = |(datain[231:228] ^ 8);
  assign w186[21] = |(datain[227:224] ^ 0);
  assign w186[22] = |(datain[223:220] ^ 15);
  assign w186[23] = |(datain[219:216] ^ 14);
  assign w186[24] = |(datain[215:212] ^ 0);
  assign w186[25] = |(datain[211:208] ^ 6);
  assign w186[26] = |(datain[207:204] ^ 7);
  assign w186[27] = |(datain[203:200] ^ 2);
  assign w186[28] = |(datain[199:196] ^ 0);
  assign w186[29] = |(datain[195:192] ^ 3);
  assign w186[30] = |(datain[191:188] ^ 14);
  assign w186[31] = |(datain[187:184] ^ 9);
  assign comp[186] = ~(|w186);
  wire [32-1:0] w187;
  assign w187[0] = |(datain[311:308] ^ 12);
  assign w187[1] = |(datain[307:304] ^ 2);
  assign w187[2] = |(datain[303:300] ^ 12);
  assign w187[3] = |(datain[299:296] ^ 5);
  assign w187[4] = |(datain[295:292] ^ 0);
  assign w187[5] = |(datain[291:288] ^ 0);
  assign w187[6] = |(datain[287:284] ^ 11);
  assign w187[7] = |(datain[283:280] ^ 4);
  assign w187[8] = |(datain[279:276] ^ 4);
  assign w187[9] = |(datain[275:272] ^ 14);
  assign w187[10] = |(datain[271:268] ^ 14);
  assign w187[11] = |(datain[267:264] ^ 11);
  assign w187[12] = |(datain[263:260] ^ 0);
  assign w187[13] = |(datain[259:256] ^ 2);
  assign w187[14] = |(datain[255:252] ^ 11);
  assign w187[15] = |(datain[251:248] ^ 4);
  assign w187[16] = |(datain[247:244] ^ 4);
  assign w187[17] = |(datain[243:240] ^ 15);
  assign w187[18] = |(datain[239:236] ^ 12);
  assign w187[19] = |(datain[235:232] ^ 13);
  assign w187[20] = |(datain[231:228] ^ 2);
  assign w187[21] = |(datain[227:224] ^ 1);
  assign w187[22] = |(datain[223:220] ^ 7);
  assign w187[23] = |(datain[219:216] ^ 3);
  assign w187[24] = |(datain[215:212] ^ 0);
  assign w187[25] = |(datain[211:208] ^ 3);
  assign w187[26] = |(datain[207:204] ^ 14);
  assign w187[27] = |(datain[203:200] ^ 9);
  assign w187[28] = |(datain[199:196] ^ 8);
  assign w187[29] = |(datain[195:192] ^ 6);
  assign w187[30] = |(datain[191:188] ^ 0);
  assign w187[31] = |(datain[187:184] ^ 0);
  assign comp[187] = ~(|w187);
  wire [42-1:0] w188;
  assign w188[0] = |(datain[311:308] ^ 0);
  assign w188[1] = |(datain[307:304] ^ 12);
  assign w188[2] = |(datain[303:300] ^ 0);
  assign w188[3] = |(datain[299:296] ^ 0);
  assign w188[4] = |(datain[295:292] ^ 11);
  assign w188[5] = |(datain[291:288] ^ 9);
  assign w188[6] = |(datain[287:284] ^ 0);
  assign w188[7] = |(datain[283:280] ^ 5);
  assign w188[8] = |(datain[279:276] ^ 0);
  assign w188[9] = |(datain[275:272] ^ 0);
  assign w188[10] = |(datain[271:268] ^ 8);
  assign w188[11] = |(datain[267:264] ^ 10);
  assign w188[12] = |(datain[263:260] ^ 0);
  assign w188[13] = |(datain[259:256] ^ 7);
  assign w188[14] = |(datain[255:252] ^ 0);
  assign w188[15] = |(datain[251:248] ^ 4);
  assign w188[16] = |(datain[247:244] ^ 1);
  assign w188[17] = |(datain[243:240] ^ 4);
  assign w188[18] = |(datain[239:236] ^ 8);
  assign w188[19] = |(datain[235:232] ^ 8);
  assign w188[20] = |(datain[231:228] ^ 4);
  assign w188[21] = |(datain[227:224] ^ 2);
  assign w188[22] = |(datain[223:220] ^ 15);
  assign w188[23] = |(datain[219:216] ^ 6);
  assign w188[24] = |(datain[215:212] ^ 4);
  assign w188[25] = |(datain[211:208] ^ 3);
  assign w188[26] = |(datain[207:204] ^ 4);
  assign w188[27] = |(datain[203:200] ^ 6);
  assign w188[28] = |(datain[199:196] ^ 14);
  assign w188[29] = |(datain[195:192] ^ 2);
  assign w188[30] = |(datain[191:188] ^ 15);
  assign w188[31] = |(datain[187:184] ^ 5);
  assign w188[32] = |(datain[183:180] ^ 12);
  assign w188[33] = |(datain[179:176] ^ 6);
  assign w188[34] = |(datain[175:172] ^ 4);
  assign w188[35] = |(datain[171:168] ^ 2);
  assign w188[36] = |(datain[167:164] ^ 15);
  assign w188[37] = |(datain[163:160] ^ 6);
  assign w188[38] = |(datain[159:156] ^ 0);
  assign w188[39] = |(datain[155:152] ^ 0);
  assign w188[40] = |(datain[151:148] ^ 12);
  assign w188[41] = |(datain[147:144] ^ 7);
  assign comp[188] = ~(|w188);
  wire [48-1:0] w189;
  assign w189[0] = |(datain[311:308] ^ 8);
  assign w189[1] = |(datain[307:304] ^ 11);
  assign w189[2] = |(datain[303:300] ^ 4);
  assign w189[3] = |(datain[299:296] ^ 6);
  assign w189[4] = |(datain[295:292] ^ 15);
  assign w189[5] = |(datain[291:288] ^ 4);
  assign w189[6] = |(datain[287:284] ^ 10);
  assign w189[7] = |(datain[283:280] ^ 3);
  assign w189[8] = |(datain[279:276] ^ 0);
  assign w189[9] = |(datain[275:272] ^ 4);
  assign w189[10] = |(datain[271:268] ^ 0);
  assign w189[11] = |(datain[267:264] ^ 0);
  assign w189[12] = |(datain[263:260] ^ 8);
  assign w189[13] = |(datain[259:256] ^ 11);
  assign w189[14] = |(datain[255:252] ^ 4);
  assign w189[15] = |(datain[251:248] ^ 6);
  assign w189[16] = |(datain[247:244] ^ 15);
  assign w189[17] = |(datain[243:240] ^ 6);
  assign w189[18] = |(datain[239:236] ^ 10);
  assign w189[19] = |(datain[235:232] ^ 3);
  assign w189[20] = |(datain[231:228] ^ 0);
  assign w189[21] = |(datain[227:224] ^ 6);
  assign w189[22] = |(datain[223:220] ^ 0);
  assign w189[23] = |(datain[219:216] ^ 0);
  assign w189[24] = |(datain[215:212] ^ 8);
  assign w189[25] = |(datain[211:208] ^ 11);
  assign w189[26] = |(datain[207:204] ^ 4);
  assign w189[27] = |(datain[203:200] ^ 6);
  assign w189[28] = |(datain[199:196] ^ 14);
  assign w189[29] = |(datain[195:192] ^ 14);
  assign w189[30] = |(datain[191:188] ^ 10);
  assign w189[31] = |(datain[187:184] ^ 3);
  assign w189[32] = |(datain[183:180] ^ 0);
  assign w189[33] = |(datain[179:176] ^ 8);
  assign w189[34] = |(datain[175:172] ^ 0);
  assign w189[35] = |(datain[171:168] ^ 0);
  assign w189[36] = |(datain[167:164] ^ 8);
  assign w189[37] = |(datain[163:160] ^ 11);
  assign w189[38] = |(datain[159:156] ^ 4);
  assign w189[39] = |(datain[155:152] ^ 6);
  assign w189[40] = |(datain[151:148] ^ 15);
  assign w189[41] = |(datain[147:144] ^ 0);
  assign w189[42] = |(datain[143:140] ^ 10);
  assign w189[43] = |(datain[139:136] ^ 3);
  assign w189[44] = |(datain[135:132] ^ 0);
  assign w189[45] = |(datain[131:128] ^ 10);
  assign w189[46] = |(datain[127:124] ^ 0);
  assign w189[47] = |(datain[123:120] ^ 0);
  assign comp[189] = ~(|w189);
  wire [32-1:0] w190;
  assign w190[0] = |(datain[311:308] ^ 8);
  assign w190[1] = |(datain[307:304] ^ 14);
  assign w190[2] = |(datain[303:300] ^ 12);
  assign w190[3] = |(datain[299:296] ^ 1);
  assign w190[4] = |(datain[295:292] ^ 0);
  assign w190[5] = |(datain[291:288] ^ 6);
  assign w190[6] = |(datain[287:284] ^ 5);
  assign w190[7] = |(datain[283:280] ^ 0);
  assign w190[8] = |(datain[279:276] ^ 11);
  assign w190[9] = |(datain[275:272] ^ 14);
  assign w190[10] = |(datain[271:268] ^ 0);
  assign w190[11] = |(datain[267:264] ^ 0);
  assign w190[12] = |(datain[263:260] ^ 0);
  assign w190[13] = |(datain[259:256] ^ 1);
  assign w190[14] = |(datain[255:252] ^ 5);
  assign w190[15] = |(datain[251:248] ^ 6);
  assign w190[16] = |(datain[247:244] ^ 3);
  assign w190[17] = |(datain[243:240] ^ 1);
  assign w190[18] = |(datain[239:236] ^ 15);
  assign w190[19] = |(datain[235:232] ^ 15);
  assign w190[20] = |(datain[231:228] ^ 11);
  assign w190[21] = |(datain[227:224] ^ 9);
  assign w190[22] = |(datain[223:220] ^ 0);
  assign w190[23] = |(datain[219:216] ^ 11);
  assign w190[24] = |(datain[215:212] ^ 0);
  assign w190[25] = |(datain[211:208] ^ 1);
  assign w190[26] = |(datain[207:204] ^ 15);
  assign w190[27] = |(datain[203:200] ^ 3);
  assign w190[28] = |(datain[199:196] ^ 10);
  assign w190[29] = |(datain[195:192] ^ 4);
  assign w190[30] = |(datain[191:188] ^ 11);
  assign w190[31] = |(datain[187:184] ^ 13);
  assign comp[190] = ~(|w190);
  wire [46-1:0] w191;
  assign w191[0] = |(datain[311:308] ^ 5);
  assign w191[1] = |(datain[307:304] ^ 1);
  assign w191[2] = |(datain[303:300] ^ 0);
  assign w191[3] = |(datain[299:296] ^ 0);
  assign w191[4] = |(datain[295:292] ^ 14);
  assign w191[5] = |(datain[291:288] ^ 11);
  assign w191[6] = |(datain[287:284] ^ 6);
  assign w191[7] = |(datain[283:280] ^ 2);
  assign w191[8] = |(datain[279:276] ^ 9);
  assign w191[9] = |(datain[275:272] ^ 0);
  assign w191[10] = |(datain[271:268] ^ 3);
  assign w191[11] = |(datain[267:264] ^ 3);
  assign w191[12] = |(datain[263:260] ^ 12);
  assign w191[13] = |(datain[259:256] ^ 0);
  assign w191[14] = |(datain[255:252] ^ 8);
  assign w191[15] = |(datain[251:248] ^ 14);
  assign w191[16] = |(datain[247:244] ^ 12);
  assign w191[17] = |(datain[243:240] ^ 0);
  assign w191[18] = |(datain[239:236] ^ 11);
  assign w191[19] = |(datain[235:232] ^ 13);
  assign w191[20] = |(datain[231:228] ^ 6);
  assign w191[21] = |(datain[227:224] ^ 12);
  assign w191[22] = |(datain[223:220] ^ 0);
  assign w191[23] = |(datain[219:216] ^ 4);
  assign w191[24] = |(datain[215:212] ^ 2);
  assign w191[25] = |(datain[211:208] ^ 6);
  assign w191[26] = |(datain[207:204] ^ 8);
  assign w191[27] = |(datain[203:200] ^ 10);
  assign w191[28] = |(datain[199:196] ^ 5);
  assign w191[29] = |(datain[195:192] ^ 6);
  assign w191[30] = |(datain[191:188] ^ 0);
  assign w191[31] = |(datain[187:184] ^ 0);
  assign w191[32] = |(datain[183:180] ^ 2);
  assign w191[33] = |(datain[179:176] ^ 14);
  assign w191[34] = |(datain[175:172] ^ 12);
  assign w191[35] = |(datain[171:168] ^ 6);
  assign w191[36] = |(datain[167:164] ^ 0);
  assign w191[37] = |(datain[163:160] ^ 6);
  assign w191[38] = |(datain[159:156] ^ 1);
  assign w191[39] = |(datain[155:152] ^ 3);
  assign w191[40] = |(datain[151:148] ^ 0);
  assign w191[41] = |(datain[147:144] ^ 5);
  assign w191[42] = |(datain[143:140] ^ 0);
  assign w191[43] = |(datain[139:136] ^ 0);
  assign w191[44] = |(datain[135:132] ^ 9);
  assign w191[45] = |(datain[131:128] ^ 0);
  assign comp[191] = ~(|w191);
  wire [42-1:0] w192;
  assign w192[0] = |(datain[311:308] ^ 2);
  assign w192[1] = |(datain[307:304] ^ 5);
  assign w192[2] = |(datain[303:300] ^ 0);
  assign w192[3] = |(datain[299:296] ^ 0);
  assign w192[4] = |(datain[295:292] ^ 15);
  assign w192[5] = |(datain[291:288] ^ 0);
  assign w192[6] = |(datain[287:284] ^ 3);
  assign w192[7] = |(datain[283:280] ^ 13);
  assign w192[8] = |(datain[279:276] ^ 0);
  assign w192[9] = |(datain[275:272] ^ 0);
  assign w192[10] = |(datain[271:268] ^ 15);
  assign w192[11] = |(datain[267:264] ^ 0);
  assign w192[12] = |(datain[263:260] ^ 7);
  assign w192[13] = |(datain[259:256] ^ 4);
  assign w192[14] = |(datain[255:252] ^ 5);
  assign w192[15] = |(datain[251:248] ^ 15);
  assign w192[16] = |(datain[247:244] ^ 8);
  assign w192[17] = |(datain[243:240] ^ 3);
  assign w192[18] = |(datain[239:236] ^ 12);
  assign w192[19] = |(datain[235:232] ^ 3);
  assign w192[20] = |(datain[231:228] ^ 1);
  assign w192[21] = |(datain[227:224] ^ 14);
  assign w192[22] = |(datain[223:220] ^ 8);
  assign w192[23] = |(datain[219:216] ^ 11);
  assign w192[24] = |(datain[215:212] ^ 13);
  assign w192[25] = |(datain[211:208] ^ 3);
  assign w192[26] = |(datain[207:204] ^ 11);
  assign w192[27] = |(datain[203:200] ^ 4);
  assign w192[28] = |(datain[199:196] ^ 3);
  assign w192[29] = |(datain[195:192] ^ 13);
  assign w192[30] = |(datain[191:188] ^ 11);
  assign w192[31] = |(datain[187:184] ^ 0);
  assign w192[32] = |(datain[183:180] ^ 0);
  assign w192[33] = |(datain[179:176] ^ 2);
  assign w192[34] = |(datain[175:172] ^ 12);
  assign w192[35] = |(datain[171:168] ^ 13);
  assign w192[36] = |(datain[167:164] ^ 2);
  assign w192[37] = |(datain[163:160] ^ 1);
  assign w192[38] = |(datain[159:156] ^ 8);
  assign w192[39] = |(datain[155:152] ^ 11);
  assign w192[40] = |(datain[151:148] ^ 13);
  assign w192[41] = |(datain[147:144] ^ 8);
  assign comp[192] = ~(|w192);
  wire [30-1:0] w193;
  assign w193[0] = |(datain[311:308] ^ 6);
  assign w193[1] = |(datain[307:304] ^ 0);
  assign w193[2] = |(datain[303:300] ^ 0);
  assign w193[3] = |(datain[299:296] ^ 1);
  assign w193[4] = |(datain[295:292] ^ 12);
  assign w193[5] = |(datain[291:288] ^ 13);
  assign w193[6] = |(datain[287:284] ^ 2);
  assign w193[7] = |(datain[283:280] ^ 1);
  assign w193[8] = |(datain[279:276] ^ 11);
  assign w193[9] = |(datain[275:272] ^ 15);
  assign w193[10] = |(datain[271:268] ^ 5);
  assign w193[11] = |(datain[267:264] ^ 2);
  assign w193[12] = |(datain[263:260] ^ 0);
  assign w193[13] = |(datain[259:256] ^ 1);
  assign w193[14] = |(datain[255:252] ^ 10);
  assign w193[15] = |(datain[251:248] ^ 1);
  assign w193[16] = |(datain[247:244] ^ 2);
  assign w193[17] = |(datain[243:240] ^ 12);
  assign w193[18] = |(datain[239:236] ^ 0);
  assign w193[19] = |(datain[235:232] ^ 0);
  assign w193[20] = |(datain[231:228] ^ 8);
  assign w193[21] = |(datain[227:224] ^ 14);
  assign w193[22] = |(datain[223:220] ^ 13);
  assign w193[23] = |(datain[219:216] ^ 8);
  assign w193[24] = |(datain[215:212] ^ 0);
  assign w193[25] = |(datain[211:208] ^ 14);
  assign w193[26] = |(datain[207:204] ^ 0);
  assign w193[27] = |(datain[203:200] ^ 7);
  assign w193[28] = |(datain[199:196] ^ 10);
  assign w193[29] = |(datain[195:192] ^ 11);
  assign comp[193] = ~(|w193);
  wire [30-1:0] w194;
  assign w194[0] = |(datain[311:308] ^ 12);
  assign w194[1] = |(datain[307:304] ^ 0);
  assign w194[2] = |(datain[303:300] ^ 0);
  assign w194[3] = |(datain[299:296] ^ 1);
  assign w194[4] = |(datain[295:292] ^ 0);
  assign w194[5] = |(datain[291:288] ^ 6);
  assign w194[6] = |(datain[287:284] ^ 14);
  assign w194[7] = |(datain[283:280] ^ 0);
  assign w194[8] = |(datain[279:276] ^ 0);
  assign w194[9] = |(datain[275:272] ^ 5);
  assign w194[10] = |(datain[271:268] ^ 0);
  assign w194[11] = |(datain[267:264] ^ 1);
  assign w194[12] = |(datain[263:260] ^ 0);
  assign w194[13] = |(datain[259:256] ^ 6);
  assign w194[14] = |(datain[255:252] ^ 4);
  assign w194[15] = |(datain[251:248] ^ 8);
  assign w194[16] = |(datain[247:244] ^ 0);
  assign w194[17] = |(datain[243:240] ^ 6);
  assign w194[18] = |(datain[239:236] ^ 10);
  assign w194[19] = |(datain[235:232] ^ 3);
  assign w194[20] = |(datain[231:228] ^ 1);
  assign w194[21] = |(datain[227:224] ^ 4);
  assign w194[22] = |(datain[223:220] ^ 0);
  assign w194[23] = |(datain[219:216] ^ 0);
  assign w194[24] = |(datain[215:212] ^ 3);
  assign w194[25] = |(datain[211:208] ^ 3);
  assign w194[26] = |(datain[207:204] ^ 12);
  assign w194[27] = |(datain[203:200] ^ 0);
  assign w194[28] = |(datain[199:196] ^ 8);
  assign w194[29] = |(datain[195:192] ^ 14);
  assign comp[194] = ~(|w194);
  wire [32-1:0] w195;
  assign w195[0] = |(datain[311:308] ^ 13);
  assign w195[1] = |(datain[307:304] ^ 2);
  assign w195[2] = |(datain[303:300] ^ 11);
  assign w195[3] = |(datain[299:296] ^ 11);
  assign w195[4] = |(datain[295:292] ^ 1);
  assign w195[5] = |(datain[291:288] ^ 0);
  assign w195[6] = |(datain[287:284] ^ 0);
  assign w195[7] = |(datain[283:280] ^ 0);
  assign w195[8] = |(datain[279:276] ^ 15);
  assign w195[9] = |(datain[275:272] ^ 7);
  assign w195[10] = |(datain[271:268] ^ 14);
  assign w195[11] = |(datain[267:264] ^ 3);
  assign w195[12] = |(datain[263:260] ^ 0);
  assign w195[13] = |(datain[259:256] ^ 3);
  assign w195[14] = |(datain[255:252] ^ 12);
  assign w195[15] = |(datain[251:248] ^ 1);
  assign w195[16] = |(datain[247:244] ^ 8);
  assign w195[17] = |(datain[243:240] ^ 3);
  assign w195[18] = |(datain[239:236] ^ 13);
  assign w195[19] = |(datain[235:232] ^ 2);
  assign w195[20] = |(datain[231:228] ^ 0);
  assign w195[21] = |(datain[227:224] ^ 0);
  assign w195[22] = |(datain[223:220] ^ 15);
  assign w195[23] = |(datain[219:216] ^ 7);
  assign w195[24] = |(datain[215:212] ^ 15);
  assign w195[25] = |(datain[211:208] ^ 3);
  assign w195[26] = |(datain[207:204] ^ 5);
  assign w195[27] = |(datain[203:200] ^ 9);
  assign w195[28] = |(datain[199:196] ^ 5);
  assign w195[29] = |(datain[195:192] ^ 0);
  assign w195[30] = |(datain[191:188] ^ 11);
  assign w195[31] = |(datain[187:184] ^ 8);
  assign comp[195] = ~(|w195);
  wire [30-1:0] w196;
  assign w196[0] = |(datain[311:308] ^ 14);
  assign w196[1] = |(datain[307:304] ^ 9);
  assign w196[2] = |(datain[303:300] ^ 1);
  assign w196[3] = |(datain[299:296] ^ 15);
  assign w196[4] = |(datain[295:292] ^ 8);
  assign w196[5] = |(datain[291:288] ^ 12);
  assign w196[6] = |(datain[287:284] ^ 12);
  assign w196[7] = |(datain[283:280] ^ 8);
  assign w196[8] = |(datain[279:276] ^ 3);
  assign w196[9] = |(datain[275:272] ^ 3);
  assign w196[10] = |(datain[271:268] ^ 13);
  assign w196[11] = |(datain[267:264] ^ 2);
  assign w196[12] = |(datain[263:260] ^ 11);
  assign w196[13] = |(datain[259:256] ^ 11);
  assign w196[14] = |(datain[255:252] ^ 1);
  assign w196[15] = |(datain[251:248] ^ 0);
  assign w196[16] = |(datain[247:244] ^ 0);
  assign w196[17] = |(datain[243:240] ^ 0);
  assign w196[18] = |(datain[239:236] ^ 15);
  assign w196[19] = |(datain[235:232] ^ 7);
  assign w196[20] = |(datain[231:228] ^ 14);
  assign w196[21] = |(datain[227:224] ^ 3);
  assign w196[22] = |(datain[223:220] ^ 0);
  assign w196[23] = |(datain[219:216] ^ 3);
  assign w196[24] = |(datain[215:212] ^ 12);
  assign w196[25] = |(datain[211:208] ^ 1);
  assign w196[26] = |(datain[207:204] ^ 8);
  assign w196[27] = |(datain[203:200] ^ 3);
  assign w196[28] = |(datain[199:196] ^ 13);
  assign w196[29] = |(datain[195:192] ^ 2);
  assign comp[196] = ~(|w196);
  wire [30-1:0] w197;
  assign w197[0] = |(datain[311:308] ^ 3);
  assign w197[1] = |(datain[307:304] ^ 5);
  assign w197[2] = |(datain[303:300] ^ 12);
  assign w197[3] = |(datain[299:296] ^ 13);
  assign w197[4] = |(datain[295:292] ^ 2);
  assign w197[5] = |(datain[291:288] ^ 1);
  assign w197[6] = |(datain[287:284] ^ 8);
  assign w197[7] = |(datain[283:280] ^ 9);
  assign w197[8] = |(datain[279:276] ^ 5);
  assign w197[9] = |(datain[275:272] ^ 14);
  assign w197[10] = |(datain[271:268] ^ 8);
  assign w197[11] = |(datain[267:264] ^ 12);
  assign w197[12] = |(datain[263:260] ^ 8);
  assign w197[13] = |(datain[259:256] ^ 12);
  assign w197[14] = |(datain[255:252] ^ 4);
  assign w197[15] = |(datain[251:248] ^ 6);
  assign w197[16] = |(datain[247:244] ^ 8);
  assign w197[17] = |(datain[243:240] ^ 14);
  assign w197[18] = |(datain[239:236] ^ 11);
  assign w197[19] = |(datain[235:232] ^ 4);
  assign w197[20] = |(datain[231:228] ^ 2);
  assign w197[21] = |(datain[227:224] ^ 5);
  assign w197[22] = |(datain[223:220] ^ 8);
  assign w197[23] = |(datain[219:216] ^ 13);
  assign w197[24] = |(datain[215:212] ^ 9);
  assign w197[25] = |(datain[211:208] ^ 4);
  assign w197[26] = |(datain[207:204] ^ 5);
  assign w197[27] = |(datain[203:200] ^ 7);
  assign w197[28] = |(datain[199:196] ^ 0);
  assign w197[29] = |(datain[195:192] ^ 1);
  assign comp[197] = ~(|w197);
  wire [46-1:0] w198;
  assign w198[0] = |(datain[311:308] ^ 5);
  assign w198[1] = |(datain[307:304] ^ 13);
  assign w198[2] = |(datain[303:300] ^ 0);
  assign w198[3] = |(datain[299:296] ^ 9);
  assign w198[4] = |(datain[295:292] ^ 12);
  assign w198[5] = |(datain[291:288] ^ 13);
  assign w198[6] = |(datain[287:284] ^ 2);
  assign w198[7] = |(datain[283:280] ^ 1);
  assign w198[8] = |(datain[279:276] ^ 11);
  assign w198[9] = |(datain[275:272] ^ 4);
  assign w198[10] = |(datain[271:268] ^ 3);
  assign w198[11] = |(datain[267:264] ^ 14);
  assign w198[12] = |(datain[263:260] ^ 12);
  assign w198[13] = |(datain[259:256] ^ 13);
  assign w198[14] = |(datain[255:252] ^ 2);
  assign w198[15] = |(datain[251:248] ^ 1);
  assign w198[16] = |(datain[247:244] ^ 11);
  assign w198[17] = |(datain[243:240] ^ 8);
  assign w198[18] = |(datain[239:236] ^ 0);
  assign w198[19] = |(datain[235:232] ^ 1);
  assign w198[20] = |(datain[231:228] ^ 4);
  assign w198[21] = |(datain[227:224] ^ 3);
  assign w198[22] = |(datain[223:220] ^ 3);
  assign w198[23] = |(datain[219:216] ^ 2);
  assign w198[24] = |(datain[215:212] ^ 14);
  assign w198[25] = |(datain[211:208] ^ 13);
  assign w198[26] = |(datain[207:204] ^ 8);
  assign w198[27] = |(datain[203:200] ^ 10);
  assign w198[28] = |(datain[199:196] ^ 4);
  assign w198[29] = |(datain[195:192] ^ 13);
  assign w198[30] = |(datain[191:188] ^ 0);
  assign w198[31] = |(datain[187:184] ^ 11);
  assign w198[32] = |(datain[183:180] ^ 12);
  assign w198[33] = |(datain[179:176] ^ 13);
  assign w198[34] = |(datain[175:172] ^ 2);
  assign w198[35] = |(datain[171:168] ^ 1);
  assign w198[36] = |(datain[167:164] ^ 12);
  assign w198[37] = |(datain[163:160] ^ 3);
  assign w198[38] = |(datain[159:156] ^ 1);
  assign w198[39] = |(datain[155:152] ^ 14);
  assign w198[40] = |(datain[151:148] ^ 0);
  assign w198[41] = |(datain[147:144] ^ 7);
  assign w198[42] = |(datain[143:140] ^ 15);
  assign w198[43] = |(datain[139:136] ^ 15);
  assign w198[44] = |(datain[135:132] ^ 14);
  assign w198[45] = |(datain[131:128] ^ 5);
  assign comp[198] = ~(|w198);
  wire [74-1:0] w199;
  assign w199[0] = |(datain[311:308] ^ 7);
  assign w199[1] = |(datain[307:304] ^ 2);
  assign w199[2] = |(datain[303:300] ^ 13);
  assign w199[3] = |(datain[299:296] ^ 12);
  assign w199[4] = |(datain[295:292] ^ 15);
  assign w199[5] = |(datain[291:288] ^ 14);
  assign w199[6] = |(datain[287:284] ^ 12);
  assign w199[7] = |(datain[283:280] ^ 4);
  assign w199[8] = |(datain[279:276] ^ 2);
  assign w199[9] = |(datain[275:272] ^ 14);
  assign w199[10] = |(datain[271:268] ^ 10);
  assign w199[11] = |(datain[267:264] ^ 3);
  assign w199[12] = |(datain[263:260] ^ 5);
  assign w199[13] = |(datain[259:256] ^ 0);
  assign w199[14] = |(datain[255:252] ^ 0);
  assign w199[15] = |(datain[251:248] ^ 1);
  assign w199[16] = |(datain[247:244] ^ 11);
  assign w199[17] = |(datain[243:240] ^ 8);
  assign w199[18] = |(datain[239:236] ^ 0);
  assign w199[19] = |(datain[235:232] ^ 0);
  assign w199[20] = |(datain[231:228] ^ 5);
  assign w199[21] = |(datain[227:224] ^ 7);
  assign w199[22] = |(datain[223:220] ^ 14);
  assign w199[23] = |(datain[219:216] ^ 8);
  assign w199[24] = |(datain[215:212] ^ 2);
  assign w199[25] = |(datain[211:208] ^ 15);
  assign w199[26] = |(datain[207:204] ^ 0);
  assign w199[27] = |(datain[203:200] ^ 0);
  assign w199[28] = |(datain[199:196] ^ 8);
  assign w199[29] = |(datain[195:192] ^ 3);
  assign w199[30] = |(datain[191:188] ^ 12);
  assign w199[31] = |(datain[187:184] ^ 9);
  assign w199[32] = |(datain[183:180] ^ 1);
  assign w199[33] = |(datain[179:176] ^ 15);
  assign w199[34] = |(datain[175:172] ^ 5);
  assign w199[35] = |(datain[171:168] ^ 1);
  assign w199[36] = |(datain[167:164] ^ 5);
  assign w199[37] = |(datain[163:160] ^ 2);
  assign w199[38] = |(datain[159:156] ^ 11);
  assign w199[39] = |(datain[155:152] ^ 4);
  assign w199[40] = |(datain[151:148] ^ 4);
  assign w199[41] = |(datain[147:144] ^ 0);
  assign w199[42] = |(datain[143:140] ^ 3);
  assign w199[43] = |(datain[139:136] ^ 3);
  assign w199[44] = |(datain[135:132] ^ 13);
  assign w199[45] = |(datain[131:128] ^ 2);
  assign w199[46] = |(datain[127:124] ^ 11);
  assign w199[47] = |(datain[123:120] ^ 9);
  assign w199[48] = |(datain[119:116] ^ 6);
  assign w199[49] = |(datain[115:112] ^ 7);
  assign w199[50] = |(datain[111:108] ^ 0);
  assign w199[51] = |(datain[107:104] ^ 1);
  assign w199[52] = |(datain[103:100] ^ 5);
  assign w199[53] = |(datain[99:96] ^ 1);
  assign w199[54] = |(datain[95:92] ^ 14);
  assign w199[55] = |(datain[91:88] ^ 8);
  assign w199[56] = |(datain[87:84] ^ 1);
  assign w199[57] = |(datain[83:80] ^ 15);
  assign w199[58] = |(datain[79:76] ^ 0);
  assign w199[59] = |(datain[75:72] ^ 0);
  assign w199[60] = |(datain[71:68] ^ 11);
  assign w199[61] = |(datain[67:64] ^ 8);
  assign w199[62] = |(datain[63:60] ^ 0);
  assign w199[63] = |(datain[59:56] ^ 0);
  assign w199[64] = |(datain[55:52] ^ 4);
  assign w199[65] = |(datain[51:48] ^ 2);
  assign w199[66] = |(datain[47:44] ^ 3);
  assign w199[67] = |(datain[43:40] ^ 3);
  assign w199[68] = |(datain[39:36] ^ 12);
  assign w199[69] = |(datain[35:32] ^ 9);
  assign w199[70] = |(datain[31:28] ^ 3);
  assign w199[71] = |(datain[27:24] ^ 3);
  assign w199[72] = |(datain[23:20] ^ 13);
  assign w199[73] = |(datain[19:16] ^ 2);
  assign comp[199] = ~(|w199);
  wire [74-1:0] w200;
  assign w200[0] = |(datain[311:308] ^ 2);
  assign w200[1] = |(datain[307:304] ^ 1);
  assign w200[2] = |(datain[303:300] ^ 11);
  assign w200[3] = |(datain[299:296] ^ 4);
  assign w200[4] = |(datain[295:292] ^ 4);
  assign w200[5] = |(datain[291:288] ^ 0);
  assign w200[6] = |(datain[287:284] ^ 8);
  assign w200[7] = |(datain[283:280] ^ 13);
  assign w200[8] = |(datain[279:276] ^ 9);
  assign w200[9] = |(datain[275:272] ^ 6);
  assign w200[10] = |(datain[271:268] ^ 0);
  assign w200[11] = |(datain[267:264] ^ 5);
  assign w200[12] = |(datain[263:260] ^ 0);
  assign w200[13] = |(datain[259:256] ^ 1);
  assign w200[14] = |(datain[255:252] ^ 11);
  assign w200[15] = |(datain[251:248] ^ 9);
  assign w200[16] = |(datain[247:244] ^ 6);
  assign w200[17] = |(datain[243:240] ^ 9);
  assign w200[18] = |(datain[239:236] ^ 0);
  assign w200[19] = |(datain[235:232] ^ 1);
  assign w200[20] = |(datain[231:228] ^ 12);
  assign w200[21] = |(datain[227:224] ^ 13);
  assign w200[22] = |(datain[223:220] ^ 2);
  assign w200[23] = |(datain[219:216] ^ 1);
  assign w200[24] = |(datain[215:212] ^ 11);
  assign w200[25] = |(datain[211:208] ^ 4);
  assign w200[26] = |(datain[207:204] ^ 3);
  assign w200[27] = |(datain[203:200] ^ 14);
  assign w200[28] = |(datain[199:196] ^ 12);
  assign w200[29] = |(datain[195:192] ^ 13);
  assign w200[30] = |(datain[191:188] ^ 2);
  assign w200[31] = |(datain[187:184] ^ 1);
  assign w200[32] = |(datain[183:180] ^ 12);
  assign w200[33] = |(datain[179:176] ^ 3);
  assign w200[34] = |(datain[175:172] ^ 12);
  assign w200[35] = |(datain[171:168] ^ 6);
  assign w200[36] = |(datain[167:164] ^ 8);
  assign w200[37] = |(datain[163:160] ^ 6);
  assign w200[38] = |(datain[159:156] ^ 5);
  assign w200[39] = |(datain[155:152] ^ 14);
  assign w200[40] = |(datain[151:148] ^ 0);
  assign w200[41] = |(datain[147:144] ^ 2);
  assign w200[42] = |(datain[143:140] ^ 0);
  assign w200[43] = |(datain[139:136] ^ 0);
  assign w200[44] = |(datain[135:132] ^ 0);
  assign w200[45] = |(datain[131:128] ^ 6);
  assign w200[46] = |(datain[127:124] ^ 11);
  assign w200[47] = |(datain[123:120] ^ 4);
  assign w200[48] = |(datain[119:116] ^ 2);
  assign w200[49] = |(datain[115:112] ^ 15);
  assign w200[50] = |(datain[111:108] ^ 12);
  assign w200[51] = |(datain[107:104] ^ 13);
  assign w200[52] = |(datain[103:100] ^ 2);
  assign w200[53] = |(datain[99:96] ^ 1);
  assign w200[54] = |(datain[95:92] ^ 0);
  assign w200[55] = |(datain[91:88] ^ 7);
  assign w200[56] = |(datain[87:84] ^ 8);
  assign w200[57] = |(datain[83:80] ^ 9);
  assign w200[58] = |(datain[79:76] ^ 9);
  assign w200[59] = |(datain[75:72] ^ 14);
  assign w200[60] = |(datain[71:68] ^ 5);
  assign w200[61] = |(datain[67:64] ^ 15);
  assign w200[62] = |(datain[63:60] ^ 0);
  assign w200[63] = |(datain[59:56] ^ 2);
  assign w200[64] = |(datain[55:52] ^ 8);
  assign w200[65] = |(datain[51:48] ^ 9);
  assign w200[66] = |(datain[47:44] ^ 9);
  assign w200[67] = |(datain[43:40] ^ 14);
  assign w200[68] = |(datain[39:36] ^ 6);
  assign w200[69] = |(datain[35:32] ^ 1);
  assign w200[70] = |(datain[31:28] ^ 0);
  assign w200[71] = |(datain[27:24] ^ 2);
  assign w200[72] = |(datain[23:20] ^ 12);
  assign w200[73] = |(datain[19:16] ^ 3);
  assign comp[200] = ~(|w200);
  wire [30-1:0] w201;
  assign w201[0] = |(datain[311:308] ^ 11);
  assign w201[1] = |(datain[307:304] ^ 15);
  assign w201[2] = |(datain[303:300] ^ 0);
  assign w201[3] = |(datain[299:296] ^ 0);
  assign w201[4] = |(datain[295:292] ^ 0);
  assign w201[5] = |(datain[291:288] ^ 1);
  assign w201[6] = |(datain[287:284] ^ 5);
  assign w201[7] = |(datain[283:280] ^ 7);
  assign w201[8] = |(datain[279:276] ^ 8);
  assign w201[9] = |(datain[275:272] ^ 11);
  assign w201[10] = |(datain[271:268] ^ 12);
  assign w201[11] = |(datain[267:264] ^ 12);
  assign w201[12] = |(datain[263:260] ^ 2);
  assign w201[13] = |(datain[259:256] ^ 11);
  assign w201[14] = |(datain[255:252] ^ 12);
  assign w201[15] = |(datain[251:248] ^ 14);
  assign w201[16] = |(datain[247:244] ^ 15);
  assign w201[17] = |(datain[243:240] ^ 3);
  assign w201[18] = |(datain[239:236] ^ 10);
  assign w201[19] = |(datain[235:232] ^ 4);
  assign w201[20] = |(datain[231:228] ^ 3);
  assign w201[21] = |(datain[227:224] ^ 3);
  assign w201[22] = |(datain[223:220] ^ 15);
  assign w201[23] = |(datain[219:216] ^ 6);
  assign w201[24] = |(datain[215:212] ^ 3);
  assign w201[25] = |(datain[211:208] ^ 3);
  assign w201[26] = |(datain[207:204] ^ 15);
  assign w201[27] = |(datain[203:200] ^ 15);
  assign w201[28] = |(datain[199:196] ^ 3);
  assign w201[29] = |(datain[195:192] ^ 3);
  assign comp[201] = ~(|w201);
  wire [32-1:0] w202;
  assign w202[0] = |(datain[311:308] ^ 11);
  assign w202[1] = |(datain[307:304] ^ 4);
  assign w202[2] = |(datain[303:300] ^ 1);
  assign w202[3] = |(datain[299:296] ^ 7);
  assign w202[4] = |(datain[295:292] ^ 8);
  assign w202[5] = |(datain[291:288] ^ 13);
  assign w202[6] = |(datain[287:284] ^ 1);
  assign w202[7] = |(datain[283:280] ^ 6);
  assign w202[8] = |(datain[279:276] ^ 5);
  assign w202[9] = |(datain[275:272] ^ 5);
  assign w202[10] = |(datain[271:268] ^ 0);
  assign w202[11] = |(datain[267:264] ^ 2);
  assign w202[12] = |(datain[263:260] ^ 12);
  assign w202[13] = |(datain[259:256] ^ 13);
  assign w202[14] = |(datain[255:252] ^ 2);
  assign w202[15] = |(datain[251:248] ^ 1);
  assign w202[16] = |(datain[247:244] ^ 11);
  assign w202[17] = |(datain[243:240] ^ 4);
  assign w202[18] = |(datain[239:236] ^ 3);
  assign w202[19] = |(datain[235:232] ^ 11);
  assign w202[20] = |(datain[231:228] ^ 8);
  assign w202[21] = |(datain[227:224] ^ 13);
  assign w202[22] = |(datain[223:220] ^ 1);
  assign w202[23] = |(datain[219:216] ^ 6);
  assign w202[24] = |(datain[215:212] ^ 7);
  assign w202[25] = |(datain[211:208] ^ 9);
  assign w202[26] = |(datain[207:204] ^ 0);
  assign w202[27] = |(datain[203:200] ^ 2);
  assign w202[28] = |(datain[199:196] ^ 12);
  assign w202[29] = |(datain[195:192] ^ 13);
  assign w202[30] = |(datain[191:188] ^ 2);
  assign w202[31] = |(datain[187:184] ^ 1);
  assign comp[202] = ~(|w202);
  wire [46-1:0] w203;
  assign w203[0] = |(datain[311:308] ^ 14);
  assign w203[1] = |(datain[307:304] ^ 8);
  assign w203[2] = |(datain[303:300] ^ 0);
  assign w203[3] = |(datain[299:296] ^ 0);
  assign w203[4] = |(datain[295:292] ^ 0);
  assign w203[5] = |(datain[291:288] ^ 0);
  assign w203[6] = |(datain[287:284] ^ 5);
  assign w203[7] = |(datain[283:280] ^ 14);
  assign w203[8] = |(datain[279:276] ^ 8);
  assign w203[9] = |(datain[275:272] ^ 3);
  assign w203[10] = |(datain[271:268] ^ 14);
  assign w203[11] = |(datain[267:264] ^ 14);
  assign w203[12] = |(datain[263:260] ^ 0);
  assign w203[13] = |(datain[259:256] ^ 4);
  assign w203[14] = |(datain[255:252] ^ 5);
  assign w203[15] = |(datain[251:248] ^ 6);
  assign w203[16] = |(datain[247:244] ^ 5);
  assign w203[17] = |(datain[243:240] ^ 0);
  assign w203[18] = |(datain[239:236] ^ 5);
  assign w203[19] = |(datain[235:232] ^ 3);
  assign w203[20] = |(datain[231:228] ^ 5);
  assign w203[21] = |(datain[227:224] ^ 1);
  assign w203[22] = |(datain[223:220] ^ 5);
  assign w203[23] = |(datain[219:216] ^ 2);
  assign w203[24] = |(datain[215:212] ^ 1);
  assign w203[25] = |(datain[211:208] ^ 14);
  assign w203[26] = |(datain[207:204] ^ 0);
  assign w203[27] = |(datain[203:200] ^ 6);
  assign w203[28] = |(datain[199:196] ^ 11);
  assign w203[29] = |(datain[195:192] ^ 4);
  assign w203[30] = |(datain[191:188] ^ 0);
  assign w203[31] = |(datain[187:184] ^ 4);
  assign w203[32] = |(datain[183:180] ^ 12);
  assign w203[33] = |(datain[179:176] ^ 13);
  assign w203[34] = |(datain[175:172] ^ 1);
  assign w203[35] = |(datain[171:168] ^ 10);
  assign w203[36] = |(datain[167:164] ^ 8);
  assign w203[37] = |(datain[163:160] ^ 0);
  assign w203[38] = |(datain[159:156] ^ 15);
  assign w203[39] = |(datain[155:152] ^ 14);
  assign w203[40] = |(datain[151:148] ^ 0);
  assign w203[41] = |(datain[147:144] ^ 8);
  assign w203[42] = |(datain[143:140] ^ 7);
  assign w203[43] = |(datain[139:136] ^ 5);
  assign w203[44] = |(datain[135:132] ^ 1);
  assign w203[45] = |(datain[131:128] ^ 2);
  assign comp[203] = ~(|w203);
  wire [74-1:0] w204;
  assign w204[0] = |(datain[311:308] ^ 8);
  assign w204[1] = |(datain[307:304] ^ 9);
  assign w204[2] = |(datain[303:300] ^ 0);
  assign w204[3] = |(datain[299:296] ^ 14);
  assign w204[4] = |(datain[295:292] ^ 11);
  assign w204[5] = |(datain[291:288] ^ 3);
  assign w204[6] = |(datain[287:284] ^ 0);
  assign w204[7] = |(datain[283:280] ^ 1);
  assign w204[8] = |(datain[279:276] ^ 11);
  assign w204[9] = |(datain[275:272] ^ 8);
  assign w204[10] = |(datain[271:268] ^ 0);
  assign w204[11] = |(datain[267:264] ^ 1);
  assign w204[12] = |(datain[263:260] ^ 0);
  assign w204[13] = |(datain[259:256] ^ 3);
  assign w204[14] = |(datain[255:252] ^ 9);
  assign w204[15] = |(datain[251:248] ^ 12);
  assign w204[16] = |(datain[247:244] ^ 2);
  assign w204[17] = |(datain[243:240] ^ 14);
  assign w204[18] = |(datain[239:236] ^ 15);
  assign w204[19] = |(datain[235:232] ^ 15);
  assign w204[20] = |(datain[231:228] ^ 1);
  assign w204[21] = |(datain[227:224] ^ 14);
  assign w204[22] = |(datain[223:220] ^ 11);
  assign w204[23] = |(datain[219:216] ^ 11);
  assign w204[24] = |(datain[215:212] ^ 0);
  assign w204[25] = |(datain[211:208] ^ 1);
  assign w204[26] = |(datain[207:204] ^ 7);
  assign w204[27] = |(datain[203:200] ^ 2);
  assign w204[28] = |(datain[199:196] ^ 1);
  assign w204[29] = |(datain[195:192] ^ 6);
  assign w204[30] = |(datain[191:188] ^ 11);
  assign w204[31] = |(datain[187:184] ^ 8);
  assign w204[32] = |(datain[183:180] ^ 0);
  assign w204[33] = |(datain[179:176] ^ 1);
  assign w204[34] = |(datain[175:172] ^ 0);
  assign w204[35] = |(datain[171:168] ^ 3);
  assign w204[36] = |(datain[167:164] ^ 5);
  assign w204[37] = |(datain[163:160] ^ 10);
  assign w204[38] = |(datain[159:156] ^ 5);
  assign w204[39] = |(datain[155:152] ^ 2);
  assign w204[40] = |(datain[151:148] ^ 11);
  assign w204[41] = |(datain[147:144] ^ 6);
  assign w204[42] = |(datain[143:140] ^ 0);
  assign w204[43] = |(datain[139:136] ^ 0);
  assign w204[44] = |(datain[135:132] ^ 11);
  assign w204[45] = |(datain[131:128] ^ 9);
  assign w204[46] = |(datain[127:124] ^ 0);
  assign w204[47] = |(datain[123:120] ^ 1);
  assign w204[48] = |(datain[119:116] ^ 0);
  assign w204[49] = |(datain[115:112] ^ 0);
  assign w204[50] = |(datain[111:108] ^ 0);
  assign w204[51] = |(datain[107:104] ^ 14);
  assign w204[52] = |(datain[103:100] ^ 0);
  assign w204[53] = |(datain[99:96] ^ 7);
  assign w204[54] = |(datain[95:92] ^ 8);
  assign w204[55] = |(datain[91:88] ^ 13);
  assign w204[56] = |(datain[87:84] ^ 1);
  assign w204[57] = |(datain[83:80] ^ 14);
  assign w204[58] = |(datain[79:76] ^ 0);
  assign w204[59] = |(datain[75:72] ^ 0);
  assign w204[60] = |(datain[71:68] ^ 0);
  assign w204[61] = |(datain[67:64] ^ 1);
  assign w204[62] = |(datain[63:60] ^ 9);
  assign w204[63] = |(datain[59:56] ^ 12);
  assign w204[64] = |(datain[55:52] ^ 2);
  assign w204[65] = |(datain[51:48] ^ 14);
  assign w204[66] = |(datain[47:44] ^ 15);
  assign w204[67] = |(datain[43:40] ^ 15);
  assign w204[68] = |(datain[39:36] ^ 1);
  assign w204[69] = |(datain[35:32] ^ 14);
  assign w204[70] = |(datain[31:28] ^ 11);
  assign w204[71] = |(datain[27:24] ^ 11);
  assign w204[72] = |(datain[23:20] ^ 0);
  assign w204[73] = |(datain[19:16] ^ 1);
  assign comp[204] = ~(|w204);
  wire [46-1:0] w205;
  assign w205[0] = |(datain[311:308] ^ 3);
  assign w205[1] = |(datain[307:304] ^ 3);
  assign w205[2] = |(datain[303:300] ^ 12);
  assign w205[3] = |(datain[299:296] ^ 0);
  assign w205[4] = |(datain[295:292] ^ 8);
  assign w205[5] = |(datain[291:288] ^ 14);
  assign w205[6] = |(datain[287:284] ^ 13);
  assign w205[7] = |(datain[283:280] ^ 8);
  assign w205[8] = |(datain[279:276] ^ 8);
  assign w205[9] = |(datain[275:272] ^ 14);
  assign w205[10] = |(datain[271:268] ^ 13);
  assign w205[11] = |(datain[267:264] ^ 0);
  assign w205[12] = |(datain[263:260] ^ 11);
  assign w205[13] = |(datain[259:256] ^ 12);
  assign w205[14] = |(datain[255:252] ^ 0);
  assign w205[15] = |(datain[251:248] ^ 0);
  assign w205[16] = |(datain[247:244] ^ 7);
  assign w205[17] = |(datain[243:240] ^ 12);
  assign w205[18] = |(datain[239:236] ^ 8);
  assign w205[19] = |(datain[235:232] ^ 11);
  assign w205[20] = |(datain[231:228] ^ 15);
  assign w205[21] = |(datain[227:224] ^ 4);
  assign w205[22] = |(datain[223:220] ^ 15);
  assign w205[23] = |(datain[219:216] ^ 11);
  assign w205[24] = |(datain[215:212] ^ 10);
  assign w205[25] = |(datain[211:208] ^ 1);
  assign w205[26] = |(datain[207:204] ^ 1);
  assign w205[27] = |(datain[203:200] ^ 3);
  assign w205[28] = |(datain[199:196] ^ 0);
  assign w205[29] = |(datain[195:192] ^ 4);
  assign w205[30] = |(datain[191:188] ^ 4);
  assign w205[31] = |(datain[187:184] ^ 8);
  assign w205[32] = |(datain[183:180] ^ 10);
  assign w205[33] = |(datain[179:176] ^ 3);
  assign w205[34] = |(datain[175:172] ^ 1);
  assign w205[35] = |(datain[171:168] ^ 3);
  assign w205[36] = |(datain[167:164] ^ 0);
  assign w205[37] = |(datain[163:160] ^ 4);
  assign w205[38] = |(datain[159:156] ^ 11);
  assign w205[39] = |(datain[155:152] ^ 1);
  assign w205[40] = |(datain[151:148] ^ 0);
  assign w205[41] = |(datain[147:144] ^ 6);
  assign w205[42] = |(datain[143:140] ^ 13);
  assign w205[43] = |(datain[139:136] ^ 3);
  assign w205[44] = |(datain[135:132] ^ 14);
  assign w205[45] = |(datain[131:128] ^ 0);
  assign comp[205] = ~(|w205);
  wire [32-1:0] w206;
  assign w206[0] = |(datain[311:308] ^ 2);
  assign w206[1] = |(datain[307:304] ^ 1);
  assign w206[2] = |(datain[303:300] ^ 3);
  assign w206[3] = |(datain[299:296] ^ 5);
  assign w206[4] = |(datain[295:292] ^ 12);
  assign w206[5] = |(datain[291:288] ^ 13);
  assign w206[6] = |(datain[287:284] ^ 2);
  assign w206[7] = |(datain[283:280] ^ 1);
  assign w206[8] = |(datain[279:276] ^ 8);
  assign w206[9] = |(datain[275:272] ^ 9);
  assign w206[10] = |(datain[271:268] ^ 1);
  assign w206[11] = |(datain[267:264] ^ 14);
  assign w206[12] = |(datain[263:260] ^ 5);
  assign w206[13] = |(datain[259:256] ^ 9);
  assign w206[14] = |(datain[255:252] ^ 0);
  assign w206[15] = |(datain[251:248] ^ 1);
  assign w206[16] = |(datain[247:244] ^ 8);
  assign w206[17] = |(datain[243:240] ^ 12);
  assign w206[18] = |(datain[239:236] ^ 0);
  assign w206[19] = |(datain[235:232] ^ 6);
  assign w206[20] = |(datain[231:228] ^ 5);
  assign w206[21] = |(datain[227:224] ^ 11);
  assign w206[22] = |(datain[223:220] ^ 0);
  assign w206[23] = |(datain[219:216] ^ 1);
  assign w206[24] = |(datain[215:212] ^ 8);
  assign w206[25] = |(datain[211:208] ^ 12);
  assign w206[26] = |(datain[207:204] ^ 12);
  assign w206[27] = |(datain[203:200] ^ 8);
  assign w206[28] = |(datain[199:196] ^ 8);
  assign w206[29] = |(datain[195:192] ^ 14);
  assign w206[30] = |(datain[191:188] ^ 13);
  assign w206[31] = |(datain[187:184] ^ 8);
  assign comp[206] = ~(|w206);
  wire [32-1:0] w207;
  assign w207[0] = |(datain[311:308] ^ 3);
  assign w207[1] = |(datain[307:304] ^ 4);
  assign w207[2] = |(datain[303:300] ^ 2);
  assign w207[3] = |(datain[299:296] ^ 14);
  assign w207[4] = |(datain[295:292] ^ 8);
  assign w207[5] = |(datain[291:288] ^ 9);
  assign w207[6] = |(datain[287:284] ^ 2);
  assign w207[7] = |(datain[283:280] ^ 6);
  assign w207[8] = |(datain[279:276] ^ 0);
  assign w207[9] = |(datain[275:272] ^ 3);
  assign w207[10] = |(datain[271:268] ^ 0);
  assign w207[11] = |(datain[267:264] ^ 1);
  assign w207[12] = |(datain[263:260] ^ 2);
  assign w207[13] = |(datain[259:256] ^ 14);
  assign w207[14] = |(datain[255:252] ^ 8);
  assign w207[15] = |(datain[251:248] ^ 12);
  assign w207[16] = |(datain[247:244] ^ 1);
  assign w207[17] = |(datain[243:240] ^ 6);
  assign w207[18] = |(datain[239:236] ^ 0);
  assign w207[19] = |(datain[235:232] ^ 5);
  assign w207[20] = |(datain[231:228] ^ 0);
  assign w207[21] = |(datain[227:224] ^ 1);
  assign w207[22] = |(datain[223:220] ^ 2);
  assign w207[23] = |(datain[219:216] ^ 14);
  assign w207[24] = |(datain[215:212] ^ 10);
  assign w207[25] = |(datain[211:208] ^ 3);
  assign w207[26] = |(datain[207:204] ^ 0);
  assign w207[27] = |(datain[203:200] ^ 7);
  assign w207[28] = |(datain[199:196] ^ 0);
  assign w207[29] = |(datain[195:192] ^ 1);
  assign w207[30] = |(datain[191:188] ^ 8);
  assign w207[31] = |(datain[187:184] ^ 13);
  assign comp[207] = ~(|w207);
  wire [28-1:0] w208;
  assign w208[0] = |(datain[311:308] ^ 4);
  assign w208[1] = |(datain[307:304] ^ 9);
  assign w208[2] = |(datain[303:300] ^ 0);
  assign w208[3] = |(datain[299:296] ^ 2);
  assign w208[4] = |(datain[295:292] ^ 2);
  assign w208[5] = |(datain[291:288] ^ 6);
  assign w208[6] = |(datain[287:284] ^ 10);
  assign w208[7] = |(datain[283:280] ^ 2);
  assign w208[8] = |(datain[279:276] ^ 4);
  assign w208[9] = |(datain[275:272] ^ 11);
  assign w208[10] = |(datain[271:268] ^ 0);
  assign w208[11] = |(datain[267:264] ^ 2);
  assign w208[12] = |(datain[263:260] ^ 2);
  assign w208[13] = |(datain[259:256] ^ 6);
  assign w208[14] = |(datain[255:252] ^ 10);
  assign w208[15] = |(datain[251:248] ^ 2);
  assign w208[16] = |(datain[247:244] ^ 8);
  assign w208[17] = |(datain[243:240] ^ 11);
  assign w208[18] = |(datain[239:236] ^ 0);
  assign w208[19] = |(datain[235:232] ^ 2);
  assign w208[20] = |(datain[231:228] ^ 5);
  assign w208[21] = |(datain[227:224] ^ 0);
  assign w208[22] = |(datain[223:220] ^ 11);
  assign w208[23] = |(datain[219:216] ^ 4);
  assign w208[24] = |(datain[215:212] ^ 1);
  assign w208[25] = |(datain[211:208] ^ 9);
  assign w208[26] = |(datain[207:204] ^ 12);
  assign w208[27] = |(datain[203:200] ^ 13);
  assign comp[208] = ~(|w208);
  wire [36-1:0] w209;
  assign w209[0] = |(datain[311:308] ^ 14);
  assign w209[1] = |(datain[307:304] ^ 12);
  assign w209[2] = |(datain[303:300] ^ 15);
  assign w209[3] = |(datain[299:296] ^ 12);
  assign w209[4] = |(datain[295:292] ^ 12);
  assign w209[5] = |(datain[291:288] ^ 3);
  assign w209[6] = |(datain[287:284] ^ 8);
  assign w209[7] = |(datain[283:280] ^ 3);
  assign w209[8] = |(datain[279:276] ^ 12);
  assign w209[9] = |(datain[275:272] ^ 3);
  assign w209[10] = |(datain[271:268] ^ 0);
  assign w209[11] = |(datain[267:264] ^ 3);
  assign w209[12] = |(datain[263:260] ^ 8);
  assign w209[13] = |(datain[259:256] ^ 1);
  assign w209[14] = |(datain[255:252] ^ 15);
  assign w209[15] = |(datain[251:248] ^ 11);
  assign w209[16] = |(datain[247:244] ^ 12);
  assign w209[17] = |(datain[243:240] ^ 12);
  assign w209[18] = |(datain[239:236] ^ 0);
  assign w209[19] = |(datain[235:232] ^ 2);
  assign w209[20] = |(datain[231:228] ^ 7);
  assign w209[21] = |(datain[227:224] ^ 2);
  assign w209[22] = |(datain[223:220] ^ 14);
  assign w209[23] = |(datain[219:216] ^ 9);
  assign w209[24] = |(datain[215:212] ^ 5);
  assign w209[25] = |(datain[211:208] ^ 11);
  assign w209[26] = |(datain[207:204] ^ 14);
  assign w209[27] = |(datain[203:200] ^ 8);
  assign w209[28] = |(datain[199:196] ^ 8);
  assign w209[29] = |(datain[195:192] ^ 9);
  assign w209[30] = |(datain[191:188] ^ 0);
  assign w209[31] = |(datain[187:184] ^ 10);
  assign w209[32] = |(datain[183:180] ^ 14);
  assign w209[33] = |(datain[179:176] ^ 4);
  assign w209[34] = |(datain[175:172] ^ 2);
  assign w209[35] = |(datain[171:168] ^ 1);
  assign comp[209] = ~(|w209);
  wire [28-1:0] w210;
  assign w210[0] = |(datain[311:308] ^ 3);
  assign w210[1] = |(datain[307:304] ^ 15);
  assign w210[2] = |(datain[303:300] ^ 12);
  assign w210[3] = |(datain[299:296] ^ 13);
  assign w210[4] = |(datain[295:292] ^ 2);
  assign w210[5] = |(datain[291:288] ^ 1);
  assign w210[6] = |(datain[287:284] ^ 2);
  assign w210[7] = |(datain[283:280] ^ 9);
  assign w210[8] = |(datain[279:276] ^ 12);
  assign w210[9] = |(datain[275:272] ^ 8);
  assign w210[10] = |(datain[271:268] ^ 5);
  assign w210[11] = |(datain[267:264] ^ 8);
  assign w210[12] = |(datain[263:260] ^ 7);
  assign w210[13] = |(datain[259:256] ^ 5);
  assign w210[14] = |(datain[255:252] ^ 13);
  assign w210[15] = |(datain[251:248] ^ 13);
  assign w210[16] = |(datain[247:244] ^ 15);
  assign w210[17] = |(datain[243:240] ^ 15);
  assign w210[18] = |(datain[239:236] ^ 14);
  assign w210[19] = |(datain[235:232] ^ 0);
  assign w210[20] = |(datain[231:228] ^ 11);
  assign w210[21] = |(datain[227:224] ^ 4);
  assign w210[22] = |(datain[223:220] ^ 4);
  assign w210[23] = |(datain[219:216] ^ 0);
  assign w210[24] = |(datain[215:212] ^ 14);
  assign w210[25] = |(datain[211:208] ^ 11);
  assign w210[26] = |(datain[207:204] ^ 15);
  assign w210[27] = |(datain[203:200] ^ 3);
  assign comp[210] = ~(|w210);
  wire [74-1:0] w211;
  assign w211[0] = |(datain[311:308] ^ 11);
  assign w211[1] = |(datain[307:304] ^ 11);
  assign w211[2] = |(datain[303:300] ^ 4);
  assign w211[3] = |(datain[299:296] ^ 0);
  assign w211[4] = |(datain[295:292] ^ 7);
  assign w211[5] = |(datain[291:288] ^ 13);
  assign w211[6] = |(datain[287:284] ^ 8);
  assign w211[7] = |(datain[283:280] ^ 10);
  assign w211[8] = |(datain[279:276] ^ 0);
  assign w211[9] = |(datain[275:272] ^ 7);
  assign w211[10] = |(datain[271:268] ^ 2);
  assign w211[11] = |(datain[267:264] ^ 4);
  assign w211[12] = |(datain[263:260] ^ 0);
  assign w211[13] = |(datain[259:256] ^ 3);
  assign w211[14] = |(datain[255:252] ^ 4);
  assign w211[15] = |(datain[251:248] ^ 0);
  assign w211[16] = |(datain[247:244] ^ 0);
  assign w211[17] = |(datain[243:240] ^ 1);
  assign w211[18] = |(datain[239:236] ^ 12);
  assign w211[19] = |(datain[235:232] ^ 0);
  assign w211[20] = |(datain[231:228] ^ 4);
  assign w211[21] = |(datain[227:224] ^ 8);
  assign w211[22] = |(datain[223:220] ^ 0);
  assign w211[23] = |(datain[219:216] ^ 1);
  assign w211[24] = |(datain[215:212] ^ 12);
  assign w211[25] = |(datain[211:208] ^ 3);
  assign w211[26] = |(datain[207:204] ^ 8);
  assign w211[27] = |(datain[203:200] ^ 11);
  assign w211[28] = |(datain[199:196] ^ 0);
  assign w211[29] = |(datain[195:192] ^ 7);
  assign w211[30] = |(datain[191:188] ^ 8);
  assign w211[31] = |(datain[187:184] ^ 14);
  assign w211[32] = |(datain[183:180] ^ 12);
  assign w211[33] = |(datain[179:176] ^ 0);
  assign w211[34] = |(datain[175:172] ^ 11);
  assign w211[35] = |(datain[171:168] ^ 14);
  assign w211[36] = |(datain[167:164] ^ 4);
  assign w211[37] = |(datain[163:160] ^ 9);
  assign w211[38] = |(datain[159:156] ^ 7);
  assign w211[39] = |(datain[155:152] ^ 13);
  assign w211[40] = |(datain[151:148] ^ 11);
  assign w211[41] = |(datain[147:144] ^ 8);
  assign w211[42] = |(datain[143:140] ^ 0);
  assign w211[43] = |(datain[139:136] ^ 5);
  assign w211[44] = |(datain[135:132] ^ 0);
  assign w211[45] = |(datain[131:128] ^ 0);
  assign w211[46] = |(datain[127:124] ^ 5);
  assign w211[47] = |(datain[123:120] ^ 0);
  assign w211[48] = |(datain[119:116] ^ 11);
  assign w211[49] = |(datain[115:112] ^ 0);
  assign w211[50] = |(datain[111:108] ^ 0);
  assign w211[51] = |(datain[107:104] ^ 0);
  assign w211[52] = |(datain[103:100] ^ 5);
  assign w211[53] = |(datain[99:96] ^ 0);
  assign w211[54] = |(datain[95:92] ^ 8);
  assign w211[55] = |(datain[91:88] ^ 9);
  assign w211[56] = |(datain[87:84] ^ 15);
  assign w211[57] = |(datain[83:80] ^ 3);
  assign w211[58] = |(datain[79:76] ^ 3);
  assign w211[59] = |(datain[75:72] ^ 1);
  assign w211[60] = |(datain[71:68] ^ 13);
  assign w211[61] = |(datain[67:64] ^ 2);
  assign w211[62] = |(datain[63:60] ^ 8);
  assign w211[63] = |(datain[59:56] ^ 10);
  assign w211[64] = |(datain[55:52] ^ 3);
  assign w211[65] = |(datain[51:48] ^ 7);
  assign w211[66] = |(datain[47:44] ^ 15);
  assign w211[67] = |(datain[43:40] ^ 14);
  assign w211[68] = |(datain[39:36] ^ 12);
  assign w211[69] = |(datain[35:32] ^ 3);
  assign w211[70] = |(datain[31:28] ^ 8);
  assign w211[71] = |(datain[27:24] ^ 11);
  assign w211[72] = |(datain[23:20] ^ 0);
  assign w211[73] = |(datain[19:16] ^ 15);
  assign comp[211] = ~(|w211);
  wire [32-1:0] w212;
  assign w212[0] = |(datain[311:308] ^ 10);
  assign w212[1] = |(datain[307:304] ^ 4);
  assign w212[2] = |(datain[303:300] ^ 8);
  assign w212[3] = |(datain[299:296] ^ 11);
  assign w212[4] = |(datain[295:292] ^ 15);
  assign w212[5] = |(datain[291:288] ^ 13);
  assign w212[6] = |(datain[287:284] ^ 12);
  assign w212[7] = |(datain[283:280] ^ 3);
  assign w212[8] = |(datain[279:276] ^ 11);
  assign w212[9] = |(datain[275:272] ^ 1);
  assign w212[10] = |(datain[271:268] ^ 0);
  assign w212[11] = |(datain[267:264] ^ 4);
  assign w212[12] = |(datain[263:260] ^ 13);
  assign w212[13] = |(datain[259:256] ^ 3);
  assign w212[14] = |(datain[255:252] ^ 14);
  assign w212[15] = |(datain[251:248] ^ 0);
  assign w212[16] = |(datain[247:244] ^ 0);
  assign w212[17] = |(datain[243:240] ^ 10);
  assign w212[18] = |(datain[239:236] ^ 12);
  assign w212[19] = |(datain[235:232] ^ 6);
  assign w212[20] = |(datain[231:228] ^ 15);
  assign w212[21] = |(datain[227:224] ^ 14);
  assign w212[22] = |(datain[223:220] ^ 12);
  assign w212[23] = |(datain[219:216] ^ 1);
  assign w212[24] = |(datain[215:212] ^ 13);
  assign w212[25] = |(datain[211:208] ^ 3);
  assign w212[26] = |(datain[207:204] ^ 14);
  assign w212[27] = |(datain[203:200] ^ 0);
  assign w212[28] = |(datain[199:196] ^ 0);
  assign w212[29] = |(datain[195:192] ^ 10);
  assign w212[30] = |(datain[191:188] ^ 12);
  assign w212[31] = |(datain[187:184] ^ 2);
  assign comp[212] = ~(|w212);
  wire [32-1:0] w213;
  assign w213[0] = |(datain[311:308] ^ 0);
  assign w213[1] = |(datain[307:304] ^ 2);
  assign w213[2] = |(datain[303:300] ^ 5);
  assign w213[3] = |(datain[299:296] ^ 6);
  assign w213[4] = |(datain[295:292] ^ 5);
  assign w213[5] = |(datain[291:288] ^ 10);
  assign w213[6] = |(datain[287:284] ^ 11);
  assign w213[7] = |(datain[283:280] ^ 9);
  assign w213[8] = |(datain[279:276] ^ 1);
  assign w213[9] = |(datain[275:272] ^ 8);
  assign w213[10] = |(datain[271:268] ^ 0);
  assign w213[11] = |(datain[267:264] ^ 0);
  assign w213[12] = |(datain[263:260] ^ 15);
  assign w213[13] = |(datain[259:256] ^ 6);
  assign w213[14] = |(datain[255:252] ^ 1);
  assign w213[15] = |(datain[251:248] ^ 4);
  assign w213[16] = |(datain[247:244] ^ 4);
  assign w213[17] = |(datain[243:240] ^ 6);
  assign w213[18] = |(datain[239:236] ^ 14);
  assign w213[19] = |(datain[235:232] ^ 2);
  assign w213[20] = |(datain[231:228] ^ 15);
  assign w213[21] = |(datain[227:224] ^ 11);
  assign w213[22] = |(datain[223:220] ^ 12);
  assign w213[23] = |(datain[219:216] ^ 13);
  assign w213[24] = |(datain[215:212] ^ 2);
  assign w213[25] = |(datain[211:208] ^ 1);
  assign w213[26] = |(datain[207:204] ^ 5);
  assign w213[27] = |(datain[203:200] ^ 14);
  assign w213[28] = |(datain[199:196] ^ 8);
  assign w213[29] = |(datain[195:192] ^ 1);
  assign w213[30] = |(datain[191:188] ^ 11);
  assign w213[31] = |(datain[187:184] ^ 12);
  assign comp[213] = ~(|w213);
  wire [30-1:0] w214;
  assign w214[0] = |(datain[311:308] ^ 0);
  assign w214[1] = |(datain[307:304] ^ 1);
  assign w214[2] = |(datain[303:300] ^ 8);
  assign w214[3] = |(datain[299:296] ^ 4);
  assign w214[4] = |(datain[295:292] ^ 10);
  assign w214[5] = |(datain[291:288] ^ 10);
  assign w214[6] = |(datain[287:284] ^ 0);
  assign w214[7] = |(datain[283:280] ^ 2);
  assign w214[8] = |(datain[279:276] ^ 2);
  assign w214[9] = |(datain[275:272] ^ 14);
  assign w214[10] = |(datain[271:268] ^ 8);
  assign w214[11] = |(datain[267:264] ^ 3);
  assign w214[12] = |(datain[263:260] ^ 8);
  assign w214[13] = |(datain[259:256] ^ 4);
  assign w214[14] = |(datain[255:252] ^ 10);
  assign w214[15] = |(datain[251:248] ^ 10);
  assign w214[16] = |(datain[247:244] ^ 0);
  assign w214[17] = |(datain[243:240] ^ 2);
  assign w214[18] = |(datain[239:236] ^ 1);
  assign w214[19] = |(datain[235:232] ^ 0);
  assign w214[20] = |(datain[231:228] ^ 0);
  assign w214[21] = |(datain[227:224] ^ 6);
  assign w214[22] = |(datain[223:220] ^ 1);
  assign w214[23] = |(datain[219:216] ^ 14);
  assign w214[24] = |(datain[215:212] ^ 11);
  assign w214[25] = |(datain[211:208] ^ 4);
  assign w214[26] = |(datain[207:204] ^ 15);
  assign w214[27] = |(datain[203:200] ^ 14);
  assign w214[28] = |(datain[199:196] ^ 12);
  assign w214[29] = |(datain[195:192] ^ 13);
  assign comp[214] = ~(|w214);
  wire [46-1:0] w215;
  assign w215[0] = |(datain[311:308] ^ 7);
  assign w215[1] = |(datain[307:304] ^ 7);
  assign w215[2] = |(datain[303:300] ^ 6);
  assign w215[3] = |(datain[299:296] ^ 7);
  assign w215[4] = |(datain[295:292] ^ 12);
  assign w215[5] = |(datain[291:288] ^ 13);
  assign w215[6] = |(datain[287:284] ^ 2);
  assign w215[7] = |(datain[283:280] ^ 1);
  assign w215[8] = |(datain[279:276] ^ 3);
  assign w215[9] = |(datain[275:272] ^ 13);
  assign w215[10] = |(datain[271:268] ^ 7);
  assign w215[11] = |(datain[267:264] ^ 3);
  assign w215[12] = |(datain[263:260] ^ 8);
  assign w215[13] = |(datain[259:256] ^ 6);
  assign w215[14] = |(datain[255:252] ^ 7);
  assign w215[15] = |(datain[251:248] ^ 4);
  assign w215[16] = |(datain[247:244] ^ 7);
  assign w215[17] = |(datain[243:240] ^ 8);
  assign w215[18] = |(datain[239:236] ^ 14);
  assign w215[19] = |(datain[235:232] ^ 8);
  assign w215[20] = |(datain[231:228] ^ 13);
  assign w215[21] = |(datain[227:224] ^ 14);
  assign w215[22] = |(datain[223:220] ^ 0);
  assign w215[23] = |(datain[219:216] ^ 3);
  assign w215[24] = |(datain[215:212] ^ 10);
  assign w215[25] = |(datain[211:208] ^ 1);
  assign w215[26] = |(datain[207:204] ^ 0);
  assign w215[27] = |(datain[203:200] ^ 15);
  assign w215[28] = |(datain[199:196] ^ 0);
  assign w215[29] = |(datain[195:192] ^ 6);
  assign w215[30] = |(datain[191:188] ^ 8);
  assign w215[31] = |(datain[187:184] ^ 0);
  assign w215[32] = |(datain[183:180] ^ 15);
  assign w215[33] = |(datain[179:176] ^ 12);
  assign w215[34] = |(datain[175:172] ^ 0);
  assign w215[35] = |(datain[171:168] ^ 4);
  assign w215[36] = |(datain[167:164] ^ 7);
  assign w215[37] = |(datain[163:160] ^ 5);
  assign w215[38] = |(datain[159:156] ^ 1);
  assign w215[39] = |(datain[155:152] ^ 0);
  assign w215[40] = |(datain[151:148] ^ 11);
  assign w215[41] = |(datain[147:144] ^ 4);
  assign w215[42] = |(datain[143:140] ^ 0);
  assign w215[43] = |(datain[139:136] ^ 0);
  assign w215[44] = |(datain[135:132] ^ 11);
  assign w215[45] = |(datain[131:128] ^ 3);
  assign comp[215] = ~(|w215);
  wire [30-1:0] w216;
  assign w216[0] = |(datain[311:308] ^ 8);
  assign w216[1] = |(datain[307:304] ^ 11);
  assign w216[2] = |(datain[303:300] ^ 13);
  assign w216[3] = |(datain[299:296] ^ 7);
  assign w216[4] = |(datain[295:292] ^ 8);
  assign w216[5] = |(datain[291:288] ^ 1);
  assign w216[6] = |(datain[287:284] ^ 12);
  assign w216[7] = |(datain[283:280] ^ 2);
  assign w216[8] = |(datain[279:276] ^ 1);
  assign w216[9] = |(datain[275:272] ^ 3);
  assign w216[10] = |(datain[271:268] ^ 0);
  assign w216[11] = |(datain[267:264] ^ 0);
  assign w216[12] = |(datain[263:260] ^ 11);
  assign w216[13] = |(datain[259:256] ^ 8);
  assign w216[14] = |(datain[255:252] ^ 0);
  assign w216[15] = |(datain[251:248] ^ 2);
  assign w216[16] = |(datain[247:244] ^ 3);
  assign w216[17] = |(datain[243:240] ^ 13);
  assign w216[18] = |(datain[239:236] ^ 12);
  assign w216[19] = |(datain[235:232] ^ 13);
  assign w216[20] = |(datain[231:228] ^ 2);
  assign w216[21] = |(datain[227:224] ^ 1);
  assign w216[22] = |(datain[223:220] ^ 7);
  assign w216[23] = |(datain[219:216] ^ 3);
  assign w216[24] = |(datain[215:212] ^ 0);
  assign w216[25] = |(datain[211:208] ^ 3);
  assign w216[26] = |(datain[207:204] ^ 14);
  assign w216[27] = |(datain[203:200] ^ 9);
  assign w216[28] = |(datain[199:196] ^ 9);
  assign w216[29] = |(datain[195:192] ^ 4);
  assign comp[216] = ~(|w216);
  wire [28-1:0] w217;
  assign w217[0] = |(datain[311:308] ^ 15);
  assign w217[1] = |(datain[307:304] ^ 3);
  assign w217[2] = |(datain[303:300] ^ 10);
  assign w217[3] = |(datain[299:296] ^ 4);
  assign w217[4] = |(datain[295:292] ^ 11);
  assign w217[5] = |(datain[291:288] ^ 8);
  assign w217[6] = |(datain[287:284] ^ 1);
  assign w217[7] = |(datain[283:280] ^ 12);
  assign w217[8] = |(datain[279:276] ^ 3);
  assign w217[9] = |(datain[275:272] ^ 5);
  assign w217[10] = |(datain[271:268] ^ 12);
  assign w217[11] = |(datain[267:264] ^ 13);
  assign w217[12] = |(datain[263:260] ^ 2);
  assign w217[13] = |(datain[259:256] ^ 1);
  assign w217[14] = |(datain[255:252] ^ 8);
  assign w217[15] = |(datain[251:248] ^ 1);
  assign w217[16] = |(datain[247:244] ^ 15);
  assign w217[17] = |(datain[243:240] ^ 11);
  assign w217[18] = |(datain[239:236] ^ 4);
  assign w217[19] = |(datain[235:232] ^ 5);
  assign w217[20] = |(datain[231:228] ^ 0);
  assign w217[21] = |(datain[227:224] ^ 2);
  assign w217[22] = |(datain[223:220] ^ 7);
  assign w217[23] = |(datain[219:216] ^ 5);
  assign w217[24] = |(datain[215:212] ^ 0);
  assign w217[25] = |(datain[211:208] ^ 8);
  assign w217[26] = |(datain[207:204] ^ 0);
  assign w217[27] = |(datain[203:200] ^ 14);
  assign comp[217] = ~(|w217);
  wire [28-1:0] w218;
  assign w218[0] = |(datain[311:308] ^ 2);
  assign w218[1] = |(datain[307:304] ^ 14);
  assign w218[2] = |(datain[303:300] ^ 10);
  assign w218[3] = |(datain[299:296] ^ 3);
  assign w218[4] = |(datain[295:292] ^ 0);
  assign w218[5] = |(datain[291:288] ^ 2);
  assign w218[6] = |(datain[287:284] ^ 0);
  assign w218[7] = |(datain[283:280] ^ 1);
  assign w218[8] = |(datain[279:276] ^ 8);
  assign w218[9] = |(datain[275:272] ^ 12);
  assign w218[10] = |(datain[271:268] ^ 1);
  assign w218[11] = |(datain[267:264] ^ 14);
  assign w218[12] = |(datain[263:260] ^ 2);
  assign w218[13] = |(datain[259:256] ^ 2);
  assign w218[14] = |(datain[255:252] ^ 0);
  assign w218[15] = |(datain[251:248] ^ 0);
  assign w218[16] = |(datain[247:244] ^ 12);
  assign w218[17] = |(datain[243:240] ^ 7);
  assign w218[18] = |(datain[239:236] ^ 0);
  assign w218[19] = |(datain[235:232] ^ 6);
  assign w218[20] = |(datain[231:228] ^ 2);
  assign w218[21] = |(datain[227:224] ^ 0);
  assign w218[22] = |(datain[223:220] ^ 0);
  assign w218[23] = |(datain[219:216] ^ 0);
  assign w218[24] = |(datain[215:212] ^ 8);
  assign w218[25] = |(datain[211:208] ^ 8);
  assign w218[26] = |(datain[207:204] ^ 0);
  assign w218[27] = |(datain[203:200] ^ 0);
  assign comp[218] = ~(|w218);
  wire [30-1:0] w219;
  assign w219[0] = |(datain[311:308] ^ 11);
  assign w219[1] = |(datain[307:304] ^ 1);
  assign w219[2] = |(datain[303:300] ^ 0);
  assign w219[3] = |(datain[299:296] ^ 4);
  assign w219[4] = |(datain[295:292] ^ 13);
  assign w219[5] = |(datain[291:288] ^ 3);
  assign w219[6] = |(datain[287:284] ^ 14);
  assign w219[7] = |(datain[283:280] ^ 8);
  assign w219[8] = |(datain[279:276] ^ 8);
  assign w219[9] = |(datain[275:272] ^ 12);
  assign w219[10] = |(datain[271:268] ^ 13);
  assign w219[11] = |(datain[267:264] ^ 11);
  assign w219[12] = |(datain[263:260] ^ 0);
  assign w219[13] = |(datain[259:256] ^ 3);
  assign w219[14] = |(datain[255:252] ^ 12);
  assign w219[15] = |(datain[251:248] ^ 3);
  assign w219[16] = |(datain[247:244] ^ 0);
  assign w219[17] = |(datain[243:240] ^ 5);
  assign w219[18] = |(datain[239:236] ^ 1);
  assign w219[19] = |(datain[235:232] ^ 0);
  assign w219[20] = |(datain[231:228] ^ 0);
  assign w219[21] = |(datain[227:224] ^ 0);
  assign w219[22] = |(datain[223:220] ^ 8);
  assign w219[23] = |(datain[219:216] ^ 14);
  assign w219[24] = |(datain[215:212] ^ 13);
  assign w219[25] = |(datain[211:208] ^ 8);
  assign w219[26] = |(datain[207:204] ^ 8);
  assign w219[27] = |(datain[203:200] ^ 12);
  assign w219[28] = |(datain[199:196] ^ 0);
  assign w219[29] = |(datain[195:192] ^ 6);
  assign comp[219] = ~(|w219);
  wire [38-1:0] w220;
  assign w220[0] = |(datain[311:308] ^ 15);
  assign w220[1] = |(datain[307:304] ^ 11);
  assign w220[2] = |(datain[303:300] ^ 10);
  assign w220[3] = |(datain[299:296] ^ 1);
  assign w220[4] = |(datain[295:292] ^ 0);
  assign w220[5] = |(datain[291:288] ^ 12);
  assign w220[6] = |(datain[287:284] ^ 0);
  assign w220[7] = |(datain[283:280] ^ 0);
  assign w220[8] = |(datain[279:276] ^ 2);
  assign w220[9] = |(datain[275:272] ^ 14);
  assign w220[10] = |(datain[271:268] ^ 10);
  assign w220[11] = |(datain[267:264] ^ 3);
  assign w220[12] = |(datain[263:260] ^ 0);
  assign w220[13] = |(datain[259:256] ^ 0);
  assign w220[14] = |(datain[255:252] ^ 0);
  assign w220[15] = |(datain[251:248] ^ 1);
  assign w220[16] = |(datain[247:244] ^ 10);
  assign w220[17] = |(datain[243:240] ^ 1);
  assign w220[18] = |(datain[239:236] ^ 0);
  assign w220[19] = |(datain[235:232] ^ 14);
  assign w220[20] = |(datain[231:228] ^ 0);
  assign w220[21] = |(datain[227:224] ^ 0);
  assign w220[22] = |(datain[223:220] ^ 2);
  assign w220[23] = |(datain[219:216] ^ 14);
  assign w220[24] = |(datain[215:212] ^ 10);
  assign w220[25] = |(datain[211:208] ^ 3);
  assign w220[26] = |(datain[207:204] ^ 0);
  assign w220[27] = |(datain[203:200] ^ 2);
  assign w220[28] = |(datain[199:196] ^ 0);
  assign w220[29] = |(datain[195:192] ^ 1);
  assign w220[30] = |(datain[191:188] ^ 8);
  assign w220[31] = |(datain[187:184] ^ 12);
  assign w220[32] = |(datain[183:180] ^ 1);
  assign w220[33] = |(datain[179:176] ^ 14);
  assign w220[34] = |(datain[175:172] ^ 2);
  assign w220[35] = |(datain[171:168] ^ 2);
  assign w220[36] = |(datain[167:164] ^ 0);
  assign w220[37] = |(datain[163:160] ^ 0);
  assign comp[220] = ~(|w220);
  wire [26-1:0] w221;
  assign w221[0] = |(datain[311:308] ^ 8);
  assign w221[1] = |(datain[307:304] ^ 14);
  assign w221[2] = |(datain[303:300] ^ 12);
  assign w221[3] = |(datain[299:296] ^ 3);
  assign w221[4] = |(datain[295:292] ^ 3);
  assign w221[5] = |(datain[291:288] ^ 11);
  assign w221[6] = |(datain[287:284] ^ 1);
  assign w221[7] = |(datain[283:280] ^ 5);
  assign w221[8] = |(datain[279:276] ^ 8);
  assign w221[9] = |(datain[275:272] ^ 14);
  assign w221[10] = |(datain[271:268] ^ 1);
  assign w221[11] = |(datain[267:264] ^ 13);
  assign w221[12] = |(datain[263:260] ^ 8);
  assign w221[13] = |(datain[259:256] ^ 11);
  assign w221[14] = |(datain[255:252] ^ 1);
  assign w221[15] = |(datain[251:248] ^ 5);
  assign w221[16] = |(datain[247:244] ^ 4);
  assign w221[17] = |(datain[243:240] ^ 10);
  assign w221[18] = |(datain[239:236] ^ 8);
  assign w221[19] = |(datain[235:232] ^ 14);
  assign w221[20] = |(datain[231:228] ^ 13);
  assign w221[21] = |(datain[227:224] ^ 10);
  assign w221[22] = |(datain[223:220] ^ 8);
  assign w221[23] = |(datain[219:216] ^ 11);
  assign w221[24] = |(datain[215:212] ^ 15);
  assign w221[25] = |(datain[211:208] ^ 1);
  assign comp[221] = ~(|w221);
  wire [30-1:0] w222;
  assign w222[0] = |(datain[311:308] ^ 5);
  assign w222[1] = |(datain[307:304] ^ 8);
  assign w222[2] = |(datain[303:300] ^ 0);
  assign w222[3] = |(datain[299:296] ^ 7);
  assign w222[4] = |(datain[295:292] ^ 2);
  assign w222[5] = |(datain[291:288] ^ 14);
  assign w222[6] = |(datain[287:284] ^ 15);
  assign w222[7] = |(datain[283:280] ^ 15);
  assign w222[8] = |(datain[279:276] ^ 2);
  assign w222[9] = |(datain[275:272] ^ 14);
  assign w222[10] = |(datain[271:268] ^ 0);
  assign w222[11] = |(datain[267:264] ^ 5);
  assign w222[12] = |(datain[263:260] ^ 0);
  assign w222[13] = |(datain[259:256] ^ 0);
  assign w222[14] = |(datain[255:252] ^ 8);
  assign w222[15] = |(datain[251:248] ^ 1);
  assign w222[16] = |(datain[247:244] ^ 3);
  assign w222[17] = |(datain[243:240] ^ 14);
  assign w222[18] = |(datain[239:236] ^ 1);
  assign w222[19] = |(datain[235:232] ^ 2);
  assign w222[20] = |(datain[231:228] ^ 0);
  assign w222[21] = |(datain[227:224] ^ 0);
  assign w222[22] = |(datain[223:220] ^ 4);
  assign w222[23] = |(datain[219:216] ^ 13);
  assign w222[24] = |(datain[215:212] ^ 5);
  assign w222[25] = |(datain[211:208] ^ 10);
  assign w222[26] = |(datain[207:204] ^ 7);
  assign w222[27] = |(datain[203:200] ^ 4);
  assign w222[28] = |(datain[199:196] ^ 0);
  assign w222[29] = |(datain[195:192] ^ 6);
  assign comp[222] = ~(|w222);
  wire [30-1:0] w223;
  assign w223[0] = |(datain[311:308] ^ 14);
  assign w223[1] = |(datain[307:304] ^ 13);
  assign w223[2] = |(datain[303:300] ^ 3);
  assign w223[3] = |(datain[299:296] ^ 1);
  assign w223[4] = |(datain[295:292] ^ 11);
  assign w223[5] = |(datain[291:288] ^ 8);
  assign w223[6] = |(datain[287:284] ^ 15);
  assign w223[7] = |(datain[283:280] ^ 1);
  assign w223[8] = |(datain[279:276] ^ 3);
  assign w223[9] = |(datain[275:272] ^ 0);
  assign w223[10] = |(datain[271:268] ^ 12);
  assign w223[11] = |(datain[267:264] ^ 13);
  assign w223[12] = |(datain[263:260] ^ 2);
  assign w223[13] = |(datain[259:256] ^ 1);
  assign w223[14] = |(datain[255:252] ^ 8);
  assign w223[15] = |(datain[251:248] ^ 12);
  assign w223[16] = |(datain[247:244] ^ 13);
  assign w223[17] = |(datain[243:240] ^ 11);
  assign w223[18] = |(datain[239:236] ^ 3);
  assign w223[19] = |(datain[235:232] ^ 12);
  assign w223[20] = |(datain[231:228] ^ 0);
  assign w223[21] = |(datain[227:224] ^ 2);
  assign w223[22] = |(datain[223:220] ^ 7);
  assign w223[23] = |(datain[219:216] ^ 2);
  assign w223[24] = |(datain[215:212] ^ 4);
  assign w223[25] = |(datain[211:208] ^ 6);
  assign w223[26] = |(datain[207:204] ^ 4);
  assign w223[27] = |(datain[203:200] ^ 11);
  assign w223[28] = |(datain[199:196] ^ 8);
  assign w223[29] = |(datain[195:192] ^ 14);
  assign comp[223] = ~(|w223);
  wire [22-1:0] w224;
  assign w224[0] = |(datain[311:308] ^ 0);
  assign w224[1] = |(datain[307:304] ^ 6);
  assign w224[2] = |(datain[303:300] ^ 0);
  assign w224[3] = |(datain[299:296] ^ 14);
  assign w224[4] = |(datain[295:292] ^ 1);
  assign w224[5] = |(datain[291:288] ^ 15);
  assign w224[6] = |(datain[287:284] ^ 1);
  assign w224[7] = |(datain[283:280] ^ 14);
  assign w224[8] = |(datain[279:276] ^ 0);
  assign w224[9] = |(datain[275:272] ^ 7);
  assign w224[10] = |(datain[271:268] ^ 11);
  assign w224[11] = |(datain[267:264] ^ 11);
  assign w224[12] = |(datain[263:260] ^ 1);
  assign w224[13] = |(datain[259:256] ^ 5);
  assign w224[14] = |(datain[255:252] ^ 0);
  assign w224[15] = |(datain[251:248] ^ 0);
  assign w224[16] = |(datain[247:244] ^ 2);
  assign w224[17] = |(datain[243:240] ^ 14);
  assign w224[18] = |(datain[239:236] ^ 8);
  assign w224[19] = |(datain[235:232] ^ 0);
  assign w224[20] = |(datain[231:228] ^ 3);
  assign w224[21] = |(datain[227:224] ^ 7);
  assign comp[224] = ~(|w224);
  wire [32-1:0] w225;
  assign w225[0] = |(datain[311:308] ^ 1);
  assign w225[1] = |(datain[307:304] ^ 15);
  assign w225[2] = |(datain[303:300] ^ 11);
  assign w225[3] = |(datain[299:296] ^ 10);
  assign w225[4] = |(datain[295:292] ^ 0);
  assign w225[5] = |(datain[291:288] ^ 0);
  assign w225[6] = |(datain[287:284] ^ 0);
  assign w225[7] = |(datain[283:280] ^ 1);
  assign w225[8] = |(datain[279:276] ^ 11);
  assign w225[9] = |(datain[275:272] ^ 9);
  assign w225[10] = |(datain[271:268] ^ 3);
  assign w225[11] = |(datain[267:264] ^ 12);
  assign w225[12] = |(datain[263:260] ^ 0);
  assign w225[13] = |(datain[259:256] ^ 2);
  assign w225[14] = |(datain[255:252] ^ 11);
  assign w225[15] = |(datain[251:248] ^ 8);
  assign w225[16] = |(datain[247:244] ^ 0);
  assign w225[17] = |(datain[243:240] ^ 0);
  assign w225[18] = |(datain[239:236] ^ 4);
  assign w225[19] = |(datain[235:232] ^ 0);
  assign w225[20] = |(datain[231:228] ^ 9);
  assign w225[21] = |(datain[227:224] ^ 12);
  assign w225[22] = |(datain[223:220] ^ 2);
  assign w225[23] = |(datain[219:216] ^ 14);
  assign w225[24] = |(datain[215:212] ^ 15);
  assign w225[25] = |(datain[211:208] ^ 15);
  assign w225[26] = |(datain[207:204] ^ 1);
  assign w225[27] = |(datain[203:200] ^ 14);
  assign w225[28] = |(datain[199:196] ^ 7);
  assign w225[29] = |(datain[195:192] ^ 13);
  assign w225[30] = |(datain[191:188] ^ 0);
  assign w225[31] = |(datain[187:184] ^ 2);
  assign comp[225] = ~(|w225);
  wire [28-1:0] w226;
  assign w226[0] = |(datain[311:308] ^ 0);
  assign w226[1] = |(datain[307:304] ^ 2);
  assign w226[2] = |(datain[303:300] ^ 3);
  assign w226[3] = |(datain[299:296] ^ 13);
  assign w226[4] = |(datain[295:292] ^ 11);
  assign w226[5] = |(datain[291:288] ^ 10);
  assign w226[6] = |(datain[287:284] ^ 1);
  assign w226[7] = |(datain[283:280] ^ 15);
  assign w226[8] = |(datain[279:276] ^ 0);
  assign w226[9] = |(datain[275:272] ^ 0);
  assign w226[10] = |(datain[271:268] ^ 0);
  assign w226[11] = |(datain[267:264] ^ 3);
  assign w226[12] = |(datain[263:260] ^ 13);
  assign w226[13] = |(datain[259:256] ^ 6);
  assign w226[14] = |(datain[255:252] ^ 12);
  assign w226[15] = |(datain[251:248] ^ 13);
  assign w226[16] = |(datain[247:244] ^ 2);
  assign w226[17] = |(datain[243:240] ^ 1);
  assign w226[18] = |(datain[239:236] ^ 7);
  assign w226[19] = |(datain[235:232] ^ 3);
  assign w226[20] = |(datain[231:228] ^ 0);
  assign w226[21] = |(datain[227:224] ^ 3);
  assign w226[22] = |(datain[223:220] ^ 14);
  assign w226[23] = |(datain[219:216] ^ 9);
  assign w226[24] = |(datain[215:212] ^ 9);
  assign w226[25] = |(datain[211:208] ^ 9);
  assign w226[26] = |(datain[207:204] ^ 0);
  assign w226[27] = |(datain[203:200] ^ 0);
  assign comp[226] = ~(|w226);
  wire [42-1:0] w227;
  assign w227[0] = |(datain[311:308] ^ 1);
  assign w227[1] = |(datain[307:304] ^ 14);
  assign w227[2] = |(datain[303:300] ^ 0);
  assign w227[3] = |(datain[299:296] ^ 6);
  assign w227[4] = |(datain[295:292] ^ 8);
  assign w227[5] = |(datain[291:288] ^ 0);
  assign w227[6] = |(datain[287:284] ^ 15);
  assign w227[7] = |(datain[283:280] ^ 12);
  assign w227[8] = |(datain[279:276] ^ 4);
  assign w227[9] = |(datain[275:272] ^ 12);
  assign w227[10] = |(datain[271:268] ^ 7);
  assign w227[11] = |(datain[267:264] ^ 4);
  assign w227[12] = |(datain[263:260] ^ 1);
  assign w227[13] = |(datain[259:256] ^ 8);
  assign w227[14] = |(datain[255:252] ^ 8);
  assign w227[15] = |(datain[251:248] ^ 0);
  assign w227[16] = |(datain[247:244] ^ 15);
  assign w227[17] = |(datain[243:240] ^ 12);
  assign w227[18] = |(datain[239:236] ^ 4);
  assign w227[19] = |(datain[235:232] ^ 11);
  assign w227[20] = |(datain[231:228] ^ 7);
  assign w227[21] = |(datain[227:224] ^ 4);
  assign w227[22] = |(datain[223:220] ^ 1);
  assign w227[23] = |(datain[219:216] ^ 3);
  assign w227[24] = |(datain[215:212] ^ 0);
  assign w227[25] = |(datain[211:208] ^ 7);
  assign w227[26] = |(datain[207:204] ^ 1);
  assign w227[27] = |(datain[203:200] ^ 15);
  assign w227[28] = |(datain[199:196] ^ 5);
  assign w227[29] = |(datain[195:192] ^ 15);
  assign w227[30] = |(datain[191:188] ^ 5);
  assign w227[31] = |(datain[187:184] ^ 14);
  assign w227[32] = |(datain[183:180] ^ 5);
  assign w227[33] = |(datain[179:176] ^ 10);
  assign w227[34] = |(datain[175:172] ^ 5);
  assign w227[35] = |(datain[171:168] ^ 9);
  assign w227[36] = |(datain[167:164] ^ 5);
  assign w227[37] = |(datain[163:160] ^ 11);
  assign w227[38] = |(datain[159:156] ^ 5);
  assign w227[39] = |(datain[155:152] ^ 8);
  assign w227[40] = |(datain[151:148] ^ 2);
  assign w227[41] = |(datain[147:144] ^ 14);
  assign comp[227] = ~(|w227);
  wire [30-1:0] w228;
  assign w228[0] = |(datain[311:308] ^ 1);
  assign w228[1] = |(datain[307:304] ^ 0);
  assign w228[2] = |(datain[303:300] ^ 0);
  assign w228[3] = |(datain[299:296] ^ 1);
  assign w228[4] = |(datain[295:292] ^ 11);
  assign w228[5] = |(datain[291:288] ^ 9);
  assign w228[6] = |(datain[287:284] ^ 3);
  assign w228[7] = |(datain[283:280] ^ 2);
  assign w228[8] = |(datain[279:276] ^ 0);
  assign w228[9] = |(datain[275:272] ^ 0);
  assign w228[10] = |(datain[271:268] ^ 8);
  assign w228[11] = |(datain[267:264] ^ 10);
  assign w228[12] = |(datain[263:260] ^ 2);
  assign w228[13] = |(datain[259:256] ^ 4);
  assign w228[14] = |(datain[255:252] ^ 8);
  assign w228[15] = |(datain[251:248] ^ 0);
  assign w228[16] = |(datain[247:244] ^ 15);
  assign w228[17] = |(datain[243:240] ^ 4);
  assign w228[18] = |(datain[239:236] ^ 13);
  assign w228[19] = |(datain[235:232] ^ 13);
  assign w228[20] = |(datain[231:228] ^ 8);
  assign w228[21] = |(datain[227:224] ^ 8);
  assign w228[22] = |(datain[223:220] ^ 2);
  assign w228[23] = |(datain[219:216] ^ 4);
  assign w228[24] = |(datain[215:212] ^ 4);
  assign w228[25] = |(datain[211:208] ^ 6);
  assign w228[26] = |(datain[207:204] ^ 14);
  assign w228[27] = |(datain[203:200] ^ 2);
  assign w228[28] = |(datain[199:196] ^ 15);
  assign w228[29] = |(datain[195:192] ^ 6);
  assign comp[228] = ~(|w228);
  wire [32-1:0] w229;
  assign w229[0] = |(datain[311:308] ^ 2);
  assign w229[1] = |(datain[307:304] ^ 4);
  assign w229[2] = |(datain[303:300] ^ 3);
  assign w229[3] = |(datain[299:296] ^ 5);
  assign w229[4] = |(datain[295:292] ^ 12);
  assign w229[5] = |(datain[291:288] ^ 13);
  assign w229[6] = |(datain[287:284] ^ 2);
  assign w229[7] = |(datain[283:280] ^ 1);
  assign w229[8] = |(datain[279:276] ^ 8);
  assign w229[9] = |(datain[275:272] ^ 9);
  assign w229[10] = |(datain[271:268] ^ 9);
  assign w229[11] = |(datain[267:264] ^ 12);
  assign w229[12] = |(datain[263:260] ^ 8);
  assign w229[13] = |(datain[259:256] ^ 15);
  assign w229[14] = |(datain[255:252] ^ 0);
  assign w229[15] = |(datain[251:248] ^ 0);
  assign w229[16] = |(datain[247:244] ^ 8);
  assign w229[17] = |(datain[243:240] ^ 12);
  assign w229[18] = |(datain[239:236] ^ 8);
  assign w229[19] = |(datain[235:232] ^ 4);
  assign w229[20] = |(datain[231:228] ^ 9);
  assign w229[21] = |(datain[227:224] ^ 1);
  assign w229[22] = |(datain[223:220] ^ 0);
  assign w229[23] = |(datain[219:216] ^ 0);
  assign w229[24] = |(datain[215:212] ^ 0);
  assign w229[25] = |(datain[211:208] ^ 7);
  assign w229[26] = |(datain[207:204] ^ 11);
  assign w229[27] = |(datain[203:200] ^ 8);
  assign w229[28] = |(datain[199:196] ^ 2);
  assign w229[29] = |(datain[195:192] ^ 4);
  assign w229[30] = |(datain[191:188] ^ 2);
  assign w229[31] = |(datain[187:184] ^ 5);
  assign comp[229] = ~(|w229);
  wire [32-1:0] w230;
  assign w230[0] = |(datain[311:308] ^ 0);
  assign w230[1] = |(datain[307:304] ^ 1);
  assign w230[2] = |(datain[303:300] ^ 4);
  assign w230[3] = |(datain[299:296] ^ 3);
  assign w230[4] = |(datain[295:292] ^ 8);
  assign w230[5] = |(datain[291:288] ^ 3);
  assign w230[6] = |(datain[287:284] ^ 14);
  assign w230[7] = |(datain[283:280] ^ 1);
  assign w230[8] = |(datain[279:276] ^ 15);
  assign w230[9] = |(datain[275:272] ^ 14);
  assign w230[10] = |(datain[271:268] ^ 11);
  assign w230[11] = |(datain[267:264] ^ 10);
  assign w230[12] = |(datain[263:260] ^ 3);
  assign w230[13] = |(datain[259:256] ^ 8);
  assign w230[14] = |(datain[255:252] ^ 0);
  assign w230[15] = |(datain[251:248] ^ 3);
  assign w230[16] = |(datain[247:244] ^ 0);
  assign w230[17] = |(datain[243:240] ^ 3);
  assign w230[18] = |(datain[239:236] ^ 13);
  assign w230[19] = |(datain[235:232] ^ 6);
  assign w230[20] = |(datain[231:228] ^ 12);
  assign w230[21] = |(datain[227:224] ^ 13);
  assign w230[22] = |(datain[223:220] ^ 2);
  assign w230[23] = |(datain[219:216] ^ 1);
  assign w230[24] = |(datain[215:212] ^ 11);
  assign w230[25] = |(datain[211:208] ^ 8);
  assign w230[26] = |(datain[207:204] ^ 0);
  assign w230[27] = |(datain[203:200] ^ 2);
  assign w230[28] = |(datain[199:196] ^ 3);
  assign w230[29] = |(datain[195:192] ^ 13);
  assign w230[30] = |(datain[191:188] ^ 11);
  assign w230[31] = |(datain[187:184] ^ 10);
  assign comp[230] = ~(|w230);
  wire [48-1:0] w231;
  assign w231[0] = |(datain[311:308] ^ 11);
  assign w231[1] = |(datain[307:304] ^ 8);
  assign w231[2] = |(datain[303:300] ^ 0);
  assign w231[3] = |(datain[299:296] ^ 0);
  assign w231[4] = |(datain[295:292] ^ 0);
  assign w231[5] = |(datain[291:288] ^ 0);
  assign w231[6] = |(datain[287:284] ^ 5);
  assign w231[7] = |(datain[283:280] ^ 0);
  assign w231[8] = |(datain[279:276] ^ 1);
  assign w231[9] = |(datain[275:272] ^ 15);
  assign w231[10] = |(datain[271:268] ^ 15);
  assign w231[11] = |(datain[267:264] ^ 10);
  assign w231[12] = |(datain[263:260] ^ 10);
  assign w231[13] = |(datain[259:256] ^ 1);
  assign w231[14] = |(datain[255:252] ^ 0);
  assign w231[15] = |(datain[251:248] ^ 4);
  assign w231[16] = |(datain[247:244] ^ 0);
  assign w231[17] = |(datain[243:240] ^ 0);
  assign w231[18] = |(datain[239:236] ^ 8);
  assign w231[19] = |(datain[235:232] ^ 9);
  assign w231[20] = |(datain[231:228] ^ 4);
  assign w231[21] = |(datain[227:224] ^ 6);
  assign w231[22] = |(datain[223:220] ^ 13);
  assign w231[23] = |(datain[219:216] ^ 12);
  assign w231[24] = |(datain[215:212] ^ 10);
  assign w231[25] = |(datain[211:208] ^ 1);
  assign w231[26] = |(datain[207:204] ^ 0);
  assign w231[27] = |(datain[203:200] ^ 6);
  assign w231[28] = |(datain[199:196] ^ 0);
  assign w231[29] = |(datain[195:192] ^ 0);
  assign w231[30] = |(datain[191:188] ^ 8);
  assign w231[31] = |(datain[187:184] ^ 9);
  assign w231[32] = |(datain[183:180] ^ 4);
  assign w231[33] = |(datain[179:176] ^ 6);
  assign w231[34] = |(datain[175:172] ^ 13);
  assign w231[35] = |(datain[171:168] ^ 14);
  assign w231[36] = |(datain[167:164] ^ 10);
  assign w231[37] = |(datain[163:160] ^ 1);
  assign w231[38] = |(datain[159:156] ^ 0);
  assign w231[39] = |(datain[155:152] ^ 12);
  assign w231[40] = |(datain[151:148] ^ 0);
  assign w231[41] = |(datain[147:144] ^ 0);
  assign w231[42] = |(datain[143:140] ^ 8);
  assign w231[43] = |(datain[139:136] ^ 9);
  assign w231[44] = |(datain[135:132] ^ 4);
  assign w231[45] = |(datain[131:128] ^ 6);
  assign w231[46] = |(datain[127:124] ^ 14);
  assign w231[47] = |(datain[123:120] ^ 0);
  assign comp[231] = ~(|w231);
  wire [50-1:0] w232;
  assign w232[0] = |(datain[311:308] ^ 11);
  assign w232[1] = |(datain[307:304] ^ 14);
  assign w232[2] = |(datain[303:300] ^ 0);
  assign w232[3] = |(datain[299:296] ^ 0);
  assign w232[4] = |(datain[295:292] ^ 0);
  assign w232[5] = |(datain[291:288] ^ 0);
  assign w232[6] = |(datain[287:284] ^ 8);
  assign w232[7] = |(datain[283:280] ^ 13);
  assign w232[8] = |(datain[279:276] ^ 8);
  assign w232[9] = |(datain[275:272] ^ 4);
  assign w232[10] = |(datain[271:268] ^ 2);
  assign w232[11] = |(datain[267:264] ^ 0);
  assign w232[12] = |(datain[263:260] ^ 0);
  assign w232[13] = |(datain[259:256] ^ 1);
  assign w232[14] = |(datain[255:252] ^ 5);
  assign w232[15] = |(datain[251:248] ^ 0);
  assign w232[16] = |(datain[247:244] ^ 8);
  assign w232[17] = |(datain[243:240] ^ 13);
  assign w232[18] = |(datain[239:236] ^ 11);
  assign w232[19] = |(datain[235:232] ^ 12);
  assign w232[20] = |(datain[231:228] ^ 2);
  assign w232[21] = |(datain[227:224] ^ 0);
  assign w232[22] = |(datain[223:220] ^ 0);
  assign w232[23] = |(datain[219:216] ^ 1);
  assign w232[24] = |(datain[215:212] ^ 11);
  assign w232[25] = |(datain[211:208] ^ 9);
  assign w232[26] = |(datain[207:204] ^ 5);
  assign w232[27] = |(datain[203:200] ^ 0);
  assign w232[28] = |(datain[199:196] ^ 0);
  assign w232[29] = |(datain[195:192] ^ 2);
  assign w232[30] = |(datain[191:188] ^ 8);
  assign w232[31] = |(datain[187:184] ^ 0);
  assign w232[32] = |(datain[183:180] ^ 0);
  assign w232[33] = |(datain[179:176] ^ 5);
  assign w232[34] = |(datain[175:172] ^ 0);
  assign w232[35] = |(datain[171:168] ^ 1);
  assign w232[36] = |(datain[167:164] ^ 4);
  assign w232[37] = |(datain[163:160] ^ 7);
  assign w232[38] = |(datain[159:156] ^ 4);
  assign w232[39] = |(datain[155:152] ^ 9);
  assign w232[40] = |(datain[151:148] ^ 7);
  assign w232[41] = |(datain[147:144] ^ 4);
  assign w232[42] = |(datain[143:140] ^ 0);
  assign w232[43] = |(datain[139:136] ^ 2);
  assign w232[44] = |(datain[135:132] ^ 14);
  assign w232[45] = |(datain[131:128] ^ 11);
  assign w232[46] = |(datain[127:124] ^ 15);
  assign w232[47] = |(datain[123:120] ^ 7);
  assign w232[48] = |(datain[119:116] ^ 12);
  assign w232[49] = |(datain[115:112] ^ 3);
  assign comp[232] = ~(|w232);
  wire [46-1:0] w233;
  assign w233[0] = |(datain[311:308] ^ 11);
  assign w233[1] = |(datain[307:304] ^ 9);
  assign w233[2] = |(datain[303:300] ^ 0);
  assign w233[3] = |(datain[299:296] ^ 0);
  assign w233[4] = |(datain[295:292] ^ 7);
  assign w233[5] = |(datain[291:288] ^ 0);
  assign w233[6] = |(datain[287:284] ^ 15);
  assign w233[7] = |(datain[283:280] ^ 2);
  assign w233[8] = |(datain[279:276] ^ 10);
  assign w233[9] = |(datain[275:272] ^ 14);
  assign w233[10] = |(datain[271:268] ^ 11);
  assign w233[11] = |(datain[267:264] ^ 9);
  assign w233[12] = |(datain[263:260] ^ 0);
  assign w233[13] = |(datain[259:256] ^ 4);
  assign w233[14] = |(datain[255:252] ^ 0);
  assign w233[15] = |(datain[251:248] ^ 0);
  assign w233[16] = |(datain[247:244] ^ 10);
  assign w233[17] = |(datain[243:240] ^ 12);
  assign w233[18] = |(datain[239:236] ^ 10);
  assign w233[19] = |(datain[235:232] ^ 14);
  assign w233[20] = |(datain[231:228] ^ 7);
  assign w233[21] = |(datain[227:224] ^ 5);
  assign w233[22] = |(datain[223:220] ^ 14);
  assign w233[23] = |(datain[219:216] ^ 14);
  assign w233[24] = |(datain[215:212] ^ 14);
  assign w233[25] = |(datain[211:208] ^ 2);
  assign w233[26] = |(datain[207:204] ^ 15);
  assign w233[27] = |(datain[203:200] ^ 10);
  assign w233[28] = |(datain[199:196] ^ 5);
  assign w233[29] = |(datain[195:192] ^ 14);
  assign w233[30] = |(datain[191:188] ^ 0);
  assign w233[31] = |(datain[187:184] ^ 7);
  assign w233[32] = |(datain[183:180] ^ 8);
  assign w233[33] = |(datain[179:176] ^ 9);
  assign w233[34] = |(datain[175:172] ^ 7);
  assign w233[35] = |(datain[171:168] ^ 12);
  assign w233[36] = |(datain[167:164] ^ 1);
  assign w233[37] = |(datain[163:160] ^ 7);
  assign w233[38] = |(datain[159:156] ^ 8);
  assign w233[39] = |(datain[155:152] ^ 9);
  assign w233[40] = |(datain[151:148] ^ 15);
  assign w233[41] = |(datain[147:144] ^ 7);
  assign w233[42] = |(datain[143:140] ^ 8);
  assign w233[43] = |(datain[139:136] ^ 3);
  assign w233[44] = |(datain[135:132] ^ 12);
  assign w233[45] = |(datain[131:128] ^ 7);
  assign comp[233] = ~(|w233);
  wire [42-1:0] w234;
  assign w234[0] = |(datain[311:308] ^ 8);
  assign w234[1] = |(datain[307:304] ^ 14);
  assign w234[2] = |(datain[303:300] ^ 13);
  assign w234[3] = |(datain[299:296] ^ 9);
  assign w234[4] = |(datain[295:292] ^ 11);
  assign w234[5] = |(datain[291:288] ^ 15);
  assign w234[6] = |(datain[287:284] ^ 15);
  assign w234[7] = |(datain[283:280] ^ 8);
  assign w234[8] = |(datain[279:276] ^ 0);
  assign w234[9] = |(datain[275:272] ^ 0);
  assign w234[10] = |(datain[271:268] ^ 10);
  assign w234[11] = |(datain[267:264] ^ 5);
  assign w234[12] = |(datain[263:260] ^ 10);
  assign w234[13] = |(datain[259:256] ^ 5);
  assign w234[14] = |(datain[255:252] ^ 11);
  assign w234[15] = |(datain[251:248] ^ 14);
  assign w234[16] = |(datain[247:244] ^ 8);
  assign w234[17] = |(datain[243:240] ^ 4);
  assign w234[18] = |(datain[239:236] ^ 0);
  assign w234[19] = |(datain[235:232] ^ 0);
  assign w234[20] = |(datain[231:228] ^ 10);
  assign w234[21] = |(datain[227:224] ^ 5);
  assign w234[22] = |(datain[223:220] ^ 10);
  assign w234[23] = |(datain[219:216] ^ 5);
  assign w234[24] = |(datain[215:212] ^ 12);
  assign w234[25] = |(datain[211:208] ^ 5);
  assign w234[26] = |(datain[207:204] ^ 4);
  assign w234[27] = |(datain[203:200] ^ 4);
  assign w234[28] = |(datain[199:196] ^ 15);
  assign w234[29] = |(datain[195:192] ^ 12);
  assign w234[30] = |(datain[191:188] ^ 0);
  assign w234[31] = |(datain[187:184] ^ 6);
  assign w234[32] = |(datain[183:180] ^ 5);
  assign w234[33] = |(datain[179:176] ^ 7);
  assign w234[34] = |(datain[175:172] ^ 11);
  assign w234[35] = |(datain[171:168] ^ 14);
  assign w234[36] = |(datain[167:164] ^ 0);
  assign w234[37] = |(datain[163:160] ^ 8);
  assign w234[38] = |(datain[159:156] ^ 0);
  assign w234[39] = |(datain[155:152] ^ 0);
  assign w234[40] = |(datain[151:148] ^ 11);
  assign w234[41] = |(datain[147:144] ^ 5);
  assign comp[234] = ~(|w234);
  wire [74-1:0] w235;
  assign w235[0] = |(datain[311:308] ^ 10);
  assign w235[1] = |(datain[307:304] ^ 6);
  assign w235[2] = |(datain[303:300] ^ 0);
  assign w235[3] = |(datain[299:296] ^ 2);
  assign w235[4] = |(datain[295:292] ^ 11);
  assign w235[5] = |(datain[291:288] ^ 10);
  assign w235[6] = |(datain[287:284] ^ 0);
  assign w235[7] = |(datain[283:280] ^ 0);
  assign w235[8] = |(datain[279:276] ^ 0);
  assign w235[9] = |(datain[275:272] ^ 0);
  assign w235[10] = |(datain[271:268] ^ 14);
  assign w235[11] = |(datain[267:264] ^ 8);
  assign w235[12] = |(datain[263:260] ^ 3);
  assign w235[13] = |(datain[259:256] ^ 12);
  assign w235[14] = |(datain[255:252] ^ 0);
  assign w235[15] = |(datain[251:248] ^ 0);
  assign w235[16] = |(datain[247:244] ^ 2);
  assign w235[17] = |(datain[243:240] ^ 14);
  assign w235[18] = |(datain[239:236] ^ 12);
  assign w235[19] = |(datain[235:232] ^ 7);
  assign w235[20] = |(datain[231:228] ^ 0);
  assign w235[21] = |(datain[227:224] ^ 6);
  assign w235[22] = |(datain[223:220] ^ 8);
  assign w235[23] = |(datain[219:216] ^ 7);
  assign w235[24] = |(datain[215:212] ^ 0);
  assign w235[25] = |(datain[211:208] ^ 1);
  assign w235[26] = |(datain[207:204] ^ 9);
  assign w235[27] = |(datain[203:200] ^ 3);
  assign w235[28] = |(datain[199:196] ^ 1);
  assign w235[29] = |(datain[195:192] ^ 9);
  assign w235[30] = |(datain[191:188] ^ 14);
  assign w235[31] = |(datain[187:184] ^ 8);
  assign w235[32] = |(datain[183:180] ^ 5);
  assign w235[33] = |(datain[179:176] ^ 11);
  assign w235[34] = |(datain[175:172] ^ 0);
  assign w235[35] = |(datain[171:168] ^ 0);
  assign w235[36] = |(datain[167:164] ^ 11);
  assign w235[37] = |(datain[163:160] ^ 4);
  assign w235[38] = |(datain[159:156] ^ 4);
  assign w235[39] = |(datain[155:152] ^ 0);
  assign w235[40] = |(datain[151:148] ^ 11);
  assign w235[41] = |(datain[147:144] ^ 9);
  assign w235[42] = |(datain[143:140] ^ 1);
  assign w235[43] = |(datain[139:136] ^ 8);
  assign w235[44] = |(datain[135:132] ^ 0);
  assign w235[45] = |(datain[131:128] ^ 0);
  assign w235[46] = |(datain[127:124] ^ 11);
  assign w235[47] = |(datain[123:120] ^ 10);
  assign w235[48] = |(datain[119:116] ^ 7);
  assign w235[49] = |(datain[115:112] ^ 5);
  assign w235[50] = |(datain[111:108] ^ 0);
  assign w235[51] = |(datain[107:104] ^ 1);
  assign w235[52] = |(datain[103:100] ^ 14);
  assign w235[53] = |(datain[99:96] ^ 8);
  assign w235[54] = |(datain[95:92] ^ 2);
  assign w235[55] = |(datain[91:88] ^ 7);
  assign w235[56] = |(datain[87:84] ^ 0);
  assign w235[57] = |(datain[83:80] ^ 0);
  assign w235[58] = |(datain[79:76] ^ 11);
  assign w235[59] = |(datain[75:72] ^ 8);
  assign w235[60] = |(datain[71:68] ^ 0);
  assign w235[61] = |(datain[67:64] ^ 1);
  assign w235[62] = |(datain[63:60] ^ 5);
  assign w235[63] = |(datain[59:56] ^ 7);
  assign w235[64] = |(datain[55:52] ^ 2);
  assign w235[65] = |(datain[51:48] ^ 14);
  assign w235[66] = |(datain[47:44] ^ 8);
  assign w235[67] = |(datain[43:40] ^ 11);
  assign w235[68] = |(datain[39:36] ^ 0);
  assign w235[69] = |(datain[35:32] ^ 14);
  assign w235[70] = |(datain[31:28] ^ 6);
  assign w235[71] = |(datain[27:24] ^ 15);
  assign w235[72] = |(datain[23:20] ^ 0);
  assign w235[73] = |(datain[19:16] ^ 1);
  assign comp[235] = ~(|w235);
  wire [28-1:0] w236;
  assign w236[0] = |(datain[311:308] ^ 7);
  assign w236[1] = |(datain[307:304] ^ 4);
  assign w236[2] = |(datain[303:300] ^ 1);
  assign w236[3] = |(datain[299:296] ^ 2);
  assign w236[4] = |(datain[295:292] ^ 8);
  assign w236[5] = |(datain[291:288] ^ 12);
  assign w236[6] = |(datain[287:284] ^ 12);
  assign w236[7] = |(datain[283:280] ^ 8);
  assign w236[8] = |(datain[279:276] ^ 11);
  assign w236[9] = |(datain[275:272] ^ 1);
  assign w236[10] = |(datain[271:268] ^ 0);
  assign w236[11] = |(datain[267:264] ^ 15);
  assign w236[12] = |(datain[263:260] ^ 13);
  assign w236[13] = |(datain[259:256] ^ 3);
  assign w236[14] = |(datain[255:252] ^ 14);
  assign w236[15] = |(datain[251:248] ^ 0);
  assign w236[16] = |(datain[247:244] ^ 3);
  assign w236[17] = |(datain[243:240] ^ 13);
  assign w236[18] = |(datain[239:236] ^ 0);
  assign w236[19] = |(datain[235:232] ^ 0);
  assign w236[20] = |(datain[231:228] ^ 8);
  assign w236[21] = |(datain[227:224] ^ 0);
  assign w236[22] = |(datain[223:220] ^ 7);
  assign w236[23] = |(datain[219:216] ^ 4);
  assign w236[24] = |(datain[215:212] ^ 0);
  assign w236[25] = |(datain[211:208] ^ 7);
  assign w236[26] = |(datain[207:204] ^ 11);
  assign w236[27] = |(datain[203:200] ^ 10);
  assign comp[236] = ~(|w236);
  wire [28-1:0] w237;
  assign w237[0] = |(datain[311:308] ^ 4);
  assign w237[1] = |(datain[307:304] ^ 5);
  assign w237[2] = |(datain[303:300] ^ 0);
  assign w237[3] = |(datain[299:296] ^ 1);
  assign w237[4] = |(datain[295:292] ^ 7);
  assign w237[5] = |(datain[291:288] ^ 5);
  assign w237[6] = |(datain[287:284] ^ 15);
  assign w237[7] = |(datain[283:280] ^ 6);
  assign w237[8] = |(datain[279:276] ^ 8);
  assign w237[9] = |(datain[275:272] ^ 3);
  assign w237[10] = |(datain[271:268] ^ 12);
  assign w237[11] = |(datain[267:264] ^ 7);
  assign w237[12] = |(datain[263:260] ^ 0);
  assign w237[13] = |(datain[259:256] ^ 4);
  assign w237[14] = |(datain[255:252] ^ 8);
  assign w237[15] = |(datain[251:248] ^ 11);
  assign w237[16] = |(datain[247:244] ^ 13);
  assign w237[17] = |(datain[243:240] ^ 7);
  assign w237[18] = |(datain[239:236] ^ 11);
  assign w237[19] = |(datain[235:232] ^ 8);
  assign w237[20] = |(datain[231:228] ^ 0);
  assign w237[21] = |(datain[227:224] ^ 2);
  assign w237[22] = |(datain[223:220] ^ 3);
  assign w237[23] = |(datain[219:216] ^ 13);
  assign w237[24] = |(datain[215:212] ^ 12);
  assign w237[25] = |(datain[211:208] ^ 13);
  assign w237[26] = |(datain[207:204] ^ 2);
  assign w237[27] = |(datain[203:200] ^ 1);
  assign comp[237] = ~(|w237);
  wire [28-1:0] w238;
  assign w238[0] = |(datain[311:308] ^ 2);
  assign w238[1] = |(datain[307:304] ^ 6);
  assign w238[2] = |(datain[303:300] ^ 8);
  assign w238[3] = |(datain[299:296] ^ 9);
  assign w238[4] = |(datain[295:292] ^ 0);
  assign w238[5] = |(datain[291:288] ^ 14);
  assign w238[6] = |(datain[287:284] ^ 3);
  assign w238[7] = |(datain[283:280] ^ 12);
  assign w238[8] = |(datain[279:276] ^ 0);
  assign w238[9] = |(datain[275:272] ^ 1);
  assign w238[10] = |(datain[271:268] ^ 12);
  assign w238[11] = |(datain[267:264] ^ 7);
  assign w238[12] = |(datain[263:260] ^ 0);
  assign w238[13] = |(datain[259:256] ^ 6);
  assign w238[14] = |(datain[255:252] ^ 8);
  assign w238[15] = |(datain[251:248] ^ 4);
  assign w238[16] = |(datain[247:244] ^ 0);
  assign w238[17] = |(datain[243:240] ^ 0);
  assign w238[18] = |(datain[239:236] ^ 2);
  assign w238[19] = |(datain[235:232] ^ 6);
  assign w238[20] = |(datain[231:228] ^ 0);
  assign w238[21] = |(datain[227:224] ^ 1);
  assign w238[22] = |(datain[223:220] ^ 8);
  assign w238[23] = |(datain[219:216] ^ 12);
  assign w238[24] = |(datain[215:212] ^ 0);
  assign w238[25] = |(datain[211:208] ^ 6);
  assign w238[26] = |(datain[207:204] ^ 8);
  assign w238[27] = |(datain[203:200] ^ 6);
  assign comp[238] = ~(|w238);
  wire [30-1:0] w239;
  assign w239[0] = |(datain[311:308] ^ 0);
  assign w239[1] = |(datain[307:304] ^ 4);
  assign w239[2] = |(datain[303:300] ^ 10);
  assign w239[3] = |(datain[299:296] ^ 1);
  assign w239[4] = |(datain[295:292] ^ 8);
  assign w239[5] = |(datain[291:288] ^ 4);
  assign w239[6] = |(datain[287:284] ^ 0);
  assign w239[7] = |(datain[283:280] ^ 0);
  assign w239[8] = |(datain[279:276] ^ 2);
  assign w239[9] = |(datain[275:272] ^ 14);
  assign w239[10] = |(datain[271:268] ^ 8);
  assign w239[11] = |(datain[267:264] ^ 9);
  assign w239[12] = |(datain[263:260] ^ 4);
  assign w239[13] = |(datain[259:256] ^ 7);
  assign w239[14] = |(datain[255:252] ^ 0);
  assign w239[15] = |(datain[251:248] ^ 11);
  assign w239[16] = |(datain[247:244] ^ 10);
  assign w239[17] = |(datain[243:240] ^ 1);
  assign w239[18] = |(datain[239:236] ^ 8);
  assign w239[19] = |(datain[235:232] ^ 6);
  assign w239[20] = |(datain[231:228] ^ 0);
  assign w239[21] = |(datain[227:224] ^ 0);
  assign w239[22] = |(datain[223:220] ^ 2);
  assign w239[23] = |(datain[219:216] ^ 14);
  assign w239[24] = |(datain[215:212] ^ 8);
  assign w239[25] = |(datain[211:208] ^ 9);
  assign w239[26] = |(datain[207:204] ^ 4);
  assign w239[27] = |(datain[203:200] ^ 7);
  assign w239[28] = |(datain[199:196] ^ 0);
  assign w239[29] = |(datain[195:192] ^ 13);
  assign comp[239] = ~(|w239);
  wire [32-1:0] w240;
  assign w240[0] = |(datain[311:308] ^ 14);
  assign w240[1] = |(datain[307:304] ^ 8);
  assign w240[2] = |(datain[303:300] ^ 10);
  assign w240[3] = |(datain[299:296] ^ 12);
  assign w240[4] = |(datain[295:292] ^ 0);
  assign w240[5] = |(datain[291:288] ^ 2);
  assign w240[6] = |(datain[287:284] ^ 14);
  assign w240[7] = |(datain[283:280] ^ 8);
  assign w240[8] = |(datain[279:276] ^ 7);
  assign w240[9] = |(datain[275:272] ^ 1);
  assign w240[10] = |(datain[271:268] ^ 0);
  assign w240[11] = |(datain[267:264] ^ 1);
  assign w240[12] = |(datain[263:260] ^ 14);
  assign w240[13] = |(datain[259:256] ^ 8);
  assign w240[14] = |(datain[255:252] ^ 9);
  assign w240[15] = |(datain[251:248] ^ 14);
  assign w240[16] = |(datain[247:244] ^ 0);
  assign w240[17] = |(datain[243:240] ^ 1);
  assign w240[18] = |(datain[239:236] ^ 14);
  assign w240[19] = |(datain[235:232] ^ 8);
  assign w240[20] = |(datain[231:228] ^ 5);
  assign w240[21] = |(datain[227:224] ^ 5);
  assign w240[22] = |(datain[223:220] ^ 0);
  assign w240[23] = |(datain[219:216] ^ 2);
  assign w240[24] = |(datain[215:212] ^ 10);
  assign w240[25] = |(datain[211:208] ^ 1);
  assign w240[26] = |(datain[207:204] ^ 2);
  assign w240[27] = |(datain[203:200] ^ 12);
  assign w240[28] = |(datain[199:196] ^ 0);
  assign w240[29] = |(datain[195:192] ^ 0);
  assign w240[30] = |(datain[191:188] ^ 8);
  assign w240[31] = |(datain[187:184] ^ 14);
  assign comp[240] = ~(|w240);
  wire [30-1:0] w241;
  assign w241[0] = |(datain[311:308] ^ 0);
  assign w241[1] = |(datain[307:304] ^ 7);
  assign w241[2] = |(datain[303:300] ^ 0);
  assign w241[3] = |(datain[299:296] ^ 0);
  assign w241[4] = |(datain[295:292] ^ 15);
  assign w241[5] = |(datain[291:288] ^ 12);
  assign w241[6] = |(datain[287:284] ^ 15);
  assign w241[7] = |(datain[283:280] ^ 3);
  assign w241[8] = |(datain[279:276] ^ 10);
  assign w241[9] = |(datain[275:272] ^ 4);
  assign w241[10] = |(datain[271:268] ^ 5);
  assign w241[11] = |(datain[267:264] ^ 8);
  assign w241[12] = |(datain[263:260] ^ 5);
  assign w241[13] = |(datain[259:256] ^ 11);
  assign w241[14] = |(datain[255:252] ^ 9);
  assign w241[15] = |(datain[251:248] ^ 13);
  assign w241[16] = |(datain[247:244] ^ 11);
  assign w241[17] = |(datain[243:240] ^ 8);
  assign w241[18] = |(datain[239:236] ^ 0);
  assign w241[19] = |(datain[235:232] ^ 0);
  assign w241[20] = |(datain[231:228] ^ 0);
  assign w241[21] = |(datain[227:224] ^ 1);
  assign w241[22] = |(datain[223:220] ^ 5);
  assign w241[23] = |(datain[219:216] ^ 3);
  assign w241[24] = |(datain[215:212] ^ 5);
  assign w241[25] = |(datain[211:208] ^ 0);
  assign w241[26] = |(datain[207:204] ^ 12);
  assign w241[27] = |(datain[203:200] ^ 11);
  assign w241[28] = |(datain[199:196] ^ 9);
  assign w241[29] = |(datain[195:192] ^ 12);
  assign comp[241] = ~(|w241);
  wire [46-1:0] w242;
  assign w242[0] = |(datain[311:308] ^ 0);
  assign w242[1] = |(datain[307:304] ^ 7);
  assign w242[2] = |(datain[303:300] ^ 0);
  assign w242[3] = |(datain[299:296] ^ 0);
  assign w242[4] = |(datain[295:292] ^ 15);
  assign w242[5] = |(datain[291:288] ^ 12);
  assign w242[6] = |(datain[287:284] ^ 15);
  assign w242[7] = |(datain[283:280] ^ 3);
  assign w242[8] = |(datain[279:276] ^ 10);
  assign w242[9] = |(datain[275:272] ^ 4);
  assign w242[10] = |(datain[271:268] ^ 5);
  assign w242[11] = |(datain[267:264] ^ 8);
  assign w242[12] = |(datain[263:260] ^ 5);
  assign w242[13] = |(datain[259:256] ^ 11);
  assign w242[14] = |(datain[255:252] ^ 9);
  assign w242[15] = |(datain[251:248] ^ 13);
  assign w242[16] = |(datain[247:244] ^ 11);
  assign w242[17] = |(datain[243:240] ^ 8);
  assign w242[18] = |(datain[239:236] ^ 0);
  assign w242[19] = |(datain[235:232] ^ 0);
  assign w242[20] = |(datain[231:228] ^ 0);
  assign w242[21] = |(datain[227:224] ^ 1);
  assign w242[22] = |(datain[223:220] ^ 5);
  assign w242[23] = |(datain[219:216] ^ 3);
  assign w242[24] = |(datain[215:212] ^ 5);
  assign w242[25] = |(datain[211:208] ^ 0);
  assign w242[26] = |(datain[207:204] ^ 12);
  assign w242[27] = |(datain[203:200] ^ 11);
  assign w242[28] = |(datain[199:196] ^ 9);
  assign w242[29] = |(datain[195:192] ^ 12);
  assign w242[30] = |(datain[191:188] ^ 3);
  assign w242[31] = |(datain[187:184] ^ 13);
  assign w242[32] = |(datain[183:180] ^ 0);
  assign w242[33] = |(datain[179:176] ^ 0);
  assign w242[34] = |(datain[175:172] ^ 12);
  assign w242[35] = |(datain[171:168] ^ 7);
  assign w242[36] = |(datain[167:164] ^ 7);
  assign w242[37] = |(datain[163:160] ^ 4);
  assign w242[38] = |(datain[159:156] ^ 13);
  assign w242[39] = |(datain[155:152] ^ 11);
  assign w242[40] = |(datain[151:148] ^ 3);
  assign w242[41] = |(datain[147:144] ^ 13);
  assign w242[42] = |(datain[143:140] ^ 0);
  assign w242[43] = |(datain[139:136] ^ 1);
  assign w242[44] = |(datain[135:132] ^ 12);
  assign w242[45] = |(datain[131:128] ^ 7);
  assign comp[242] = ~(|w242);
  wire [44-1:0] w243;
  assign w243[0] = |(datain[311:308] ^ 3);
  assign w243[1] = |(datain[307:304] ^ 6);
  assign w243[2] = |(datain[303:300] ^ 8);
  assign w243[3] = |(datain[299:296] ^ 14);
  assign w243[4] = |(datain[295:292] ^ 4);
  assign w243[5] = |(datain[291:288] ^ 6);
  assign w243[6] = |(datain[287:284] ^ 0);
  assign w243[7] = |(datain[283:280] ^ 2);
  assign w243[8] = |(datain[279:276] ^ 8);
  assign w243[9] = |(datain[275:272] ^ 11);
  assign w243[10] = |(datain[271:268] ^ 7);
  assign w243[11] = |(datain[267:264] ^ 6);
  assign w243[12] = |(datain[263:260] ^ 0);
  assign w243[13] = |(datain[259:256] ^ 10);
  assign w243[14] = |(datain[255:252] ^ 2);
  assign w243[15] = |(datain[251:248] ^ 6);
  assign w243[16] = |(datain[247:244] ^ 8);
  assign w243[17] = |(datain[243:240] ^ 10);
  assign w243[18] = |(datain[239:236] ^ 1);
  assign w243[19] = |(datain[235:232] ^ 4);
  assign w243[20] = |(datain[231:228] ^ 8);
  assign w243[21] = |(datain[227:224] ^ 0);
  assign w243[22] = |(datain[223:220] ^ 14);
  assign w243[23] = |(datain[219:216] ^ 10);
  assign w243[24] = |(datain[215:212] ^ 4);
  assign w243[25] = |(datain[211:208] ^ 0);
  assign w243[26] = |(datain[207:204] ^ 12);
  assign w243[27] = |(datain[203:200] ^ 13);
  assign w243[28] = |(datain[199:196] ^ 2);
  assign w243[29] = |(datain[195:192] ^ 1);
  assign w243[30] = |(datain[191:188] ^ 3);
  assign w243[31] = |(datain[187:184] ^ 13);
  assign w243[32] = |(datain[183:180] ^ 15);
  assign w243[33] = |(datain[179:176] ^ 15);
  assign w243[34] = |(datain[175:172] ^ 15);
  assign w243[35] = |(datain[171:168] ^ 15);
  assign w243[36] = |(datain[167:164] ^ 7);
  assign w243[37] = |(datain[163:160] ^ 4);
  assign w243[38] = |(datain[159:156] ^ 0);
  assign w243[39] = |(datain[155:152] ^ 14);
  assign w243[40] = |(datain[151:148] ^ 15);
  assign w243[41] = |(datain[147:144] ^ 7);
  assign w243[42] = |(datain[143:140] ^ 14);
  assign w243[43] = |(datain[139:136] ^ 3);
  assign comp[243] = ~(|w243);
  wire [28-1:0] w244;
  assign w244[0] = |(datain[311:308] ^ 0);
  assign w244[1] = |(datain[307:304] ^ 10);
  assign w244[2] = |(datain[303:300] ^ 2);
  assign w244[3] = |(datain[299:296] ^ 6);
  assign w244[4] = |(datain[295:292] ^ 8);
  assign w244[5] = |(datain[291:288] ^ 10);
  assign w244[6] = |(datain[287:284] ^ 1);
  assign w244[7] = |(datain[283:280] ^ 4);
  assign w244[8] = |(datain[279:276] ^ 8);
  assign w244[9] = |(datain[275:272] ^ 0);
  assign w244[10] = |(datain[271:268] ^ 14);
  assign w244[11] = |(datain[267:264] ^ 10);
  assign w244[12] = |(datain[263:260] ^ 4);
  assign w244[13] = |(datain[259:256] ^ 0);
  assign w244[14] = |(datain[255:252] ^ 12);
  assign w244[15] = |(datain[251:248] ^ 13);
  assign w244[16] = |(datain[247:244] ^ 2);
  assign w244[17] = |(datain[243:240] ^ 1);
  assign w244[18] = |(datain[239:236] ^ 3);
  assign w244[19] = |(datain[235:232] ^ 13);
  assign w244[20] = |(datain[231:228] ^ 15);
  assign w244[21] = |(datain[227:224] ^ 15);
  assign w244[22] = |(datain[223:220] ^ 15);
  assign w244[23] = |(datain[219:216] ^ 15);
  assign w244[24] = |(datain[215:212] ^ 7);
  assign w244[25] = |(datain[211:208] ^ 4);
  assign w244[26] = |(datain[207:204] ^ 0);
  assign w244[27] = |(datain[203:200] ^ 14);
  assign comp[244] = ~(|w244);
  wire [42-1:0] w245;
  assign w245[0] = |(datain[311:308] ^ 1);
  assign w245[1] = |(datain[307:304] ^ 14);
  assign w245[2] = |(datain[303:300] ^ 5);
  assign w245[3] = |(datain[299:296] ^ 7);
  assign w245[4] = |(datain[295:292] ^ 14);
  assign w245[5] = |(datain[291:288] ^ 8);
  assign w245[6] = |(datain[287:284] ^ 1);
  assign w245[7] = |(datain[283:280] ^ 8);
  assign w245[8] = |(datain[279:276] ^ 15);
  assign w245[9] = |(datain[275:272] ^ 14);
  assign w245[10] = |(datain[271:268] ^ 0);
  assign w245[11] = |(datain[267:264] ^ 8);
  assign w245[12] = |(datain[263:260] ^ 12);
  assign w245[13] = |(datain[259:256] ^ 0);
  assign w245[14] = |(datain[255:252] ^ 7);
  assign w245[15] = |(datain[251:248] ^ 4);
  assign w245[16] = |(datain[247:244] ^ 0);
  assign w245[17] = |(datain[243:240] ^ 3);
  assign w245[18] = |(datain[239:236] ^ 14);
  assign w245[19] = |(datain[235:232] ^ 9);
  assign w245[20] = |(datain[231:228] ^ 15);
  assign w245[21] = |(datain[227:224] ^ 14);
  assign w245[22] = |(datain[223:220] ^ 0);
  assign w245[23] = |(datain[219:216] ^ 0);
  assign w245[24] = |(datain[215:212] ^ 8);
  assign w245[25] = |(datain[211:208] ^ 0);
  assign w245[26] = |(datain[207:204] ^ 3);
  assign w245[27] = |(datain[203:200] ^ 14);
  assign w245[28] = |(datain[199:196] ^ 4);
  assign w245[29] = |(datain[195:192] ^ 1);
  assign w245[30] = |(datain[191:188] ^ 0);
  assign w245[31] = |(datain[187:184] ^ 0);
  assign w245[32] = |(datain[183:180] ^ 4);
  assign w245[33] = |(datain[179:176] ^ 3);
  assign w245[34] = |(datain[175:172] ^ 7);
  assign w245[35] = |(datain[171:168] ^ 5);
  assign w245[36] = |(datain[167:164] ^ 2);
  assign w245[37] = |(datain[163:160] ^ 13);
  assign w245[38] = |(datain[159:156] ^ 8);
  assign w245[39] = |(datain[155:152] ^ 0);
  assign w245[40] = |(datain[151:148] ^ 3);
  assign w245[41] = |(datain[147:144] ^ 14);
  assign comp[245] = ~(|w245);
  wire [30-1:0] w246;
  assign w246[0] = |(datain[311:308] ^ 12);
  assign w246[1] = |(datain[307:304] ^ 10);
  assign w246[2] = |(datain[303:300] ^ 0);
  assign w246[3] = |(datain[299:296] ^ 0);
  assign w246[4] = |(datain[295:292] ^ 8);
  assign w246[5] = |(datain[291:288] ^ 0);
  assign w246[6] = |(datain[287:284] ^ 3);
  assign w246[7] = |(datain[283:280] ^ 14);
  assign w246[8] = |(datain[279:276] ^ 6);
  assign w246[9] = |(datain[275:272] ^ 12);
  assign w246[10] = |(datain[271:268] ^ 4);
  assign w246[11] = |(datain[267:264] ^ 6);
  assign w246[12] = |(datain[263:260] ^ 0);
  assign w246[13] = |(datain[259:256] ^ 0);
  assign w246[14] = |(datain[255:252] ^ 7);
  assign w246[15] = |(datain[251:248] ^ 4);
  assign w246[16] = |(datain[247:244] ^ 0);
  assign w246[17] = |(datain[243:240] ^ 3);
  assign w246[18] = |(datain[239:236] ^ 14);
  assign w246[19] = |(datain[235:232] ^ 9);
  assign w246[20] = |(datain[231:228] ^ 12);
  assign w246[21] = |(datain[227:224] ^ 0);
  assign w246[22] = |(datain[223:220] ^ 0);
  assign w246[23] = |(datain[219:216] ^ 0);
  assign w246[24] = |(datain[215:212] ^ 11);
  assign w246[25] = |(datain[211:208] ^ 15);
  assign w246[26] = |(datain[207:204] ^ 14);
  assign w246[27] = |(datain[203:200] ^ 10);
  assign w246[28] = |(datain[199:196] ^ 4);
  assign w246[29] = |(datain[195:192] ^ 2);
  assign comp[246] = ~(|w246);
  wire [30-1:0] w247;
  assign w247[0] = |(datain[311:308] ^ 13);
  assign w247[1] = |(datain[307:304] ^ 5);
  assign w247[2] = |(datain[303:300] ^ 10);
  assign w247[3] = |(datain[299:296] ^ 1);
  assign w247[4] = |(datain[295:292] ^ 12);
  assign w247[5] = |(datain[291:288] ^ 13);
  assign w247[6] = |(datain[287:284] ^ 2);
  assign w247[7] = |(datain[283:280] ^ 1);
  assign w247[8] = |(datain[279:276] ^ 3);
  assign w247[9] = |(datain[275:272] ^ 13);
  assign w247[10] = |(datain[271:268] ^ 0);
  assign w247[11] = |(datain[267:264] ^ 13);
  assign w247[12] = |(datain[263:260] ^ 9);
  assign w247[13] = |(datain[259:256] ^ 0);
  assign w247[14] = |(datain[255:252] ^ 7);
  assign w247[15] = |(datain[251:248] ^ 4);
  assign w247[16] = |(datain[247:244] ^ 0);
  assign w247[17] = |(datain[243:240] ^ 9);
  assign w247[18] = |(datain[239:236] ^ 11);
  assign w247[19] = |(datain[235:232] ^ 4);
  assign w247[20] = |(datain[231:228] ^ 4);
  assign w247[21] = |(datain[227:224] ^ 10);
  assign w247[22] = |(datain[223:220] ^ 11);
  assign w247[23] = |(datain[219:216] ^ 11);
  assign w247[24] = |(datain[215:212] ^ 0);
  assign w247[25] = |(datain[211:208] ^ 0);
  assign w247[26] = |(datain[207:204] ^ 1);
  assign w247[27] = |(datain[203:200] ^ 0);
  assign w247[28] = |(datain[199:196] ^ 12);
  assign w247[29] = |(datain[195:192] ^ 13);
  assign comp[247] = ~(|w247);
  wire [24-1:0] w248;
  assign w248[0] = |(datain[311:308] ^ 13);
  assign w248[1] = |(datain[307:304] ^ 5);
  assign w248[2] = |(datain[303:300] ^ 10);
  assign w248[3] = |(datain[299:296] ^ 1);
  assign w248[4] = |(datain[295:292] ^ 7);
  assign w248[5] = |(datain[291:288] ^ 5);
  assign w248[6] = |(datain[287:284] ^ 0);
  assign w248[7] = |(datain[283:280] ^ 5);
  assign w248[8] = |(datain[279:276] ^ 11);
  assign w248[9] = |(datain[275:272] ^ 8);
  assign w248[10] = |(datain[271:268] ^ 0);
  assign w248[11] = |(datain[267:264] ^ 13);
  assign w248[12] = |(datain[263:260] ^ 9);
  assign w248[13] = |(datain[259:256] ^ 0);
  assign w248[14] = |(datain[255:252] ^ 9);
  assign w248[15] = |(datain[251:248] ^ 13);
  assign w248[16] = |(datain[247:244] ^ 12);
  assign w248[17] = |(datain[243:240] ^ 15);
  assign w248[18] = |(datain[239:236] ^ 2);
  assign w248[19] = |(datain[235:232] ^ 14);
  assign w248[20] = |(datain[231:228] ^ 15);
  assign w248[21] = |(datain[227:224] ^ 15);
  assign w248[22] = |(datain[223:220] ^ 3);
  assign w248[23] = |(datain[219:216] ^ 6);
  assign comp[248] = ~(|w248);
  wire [76-1:0] w249;
  assign w249[0] = |(datain[311:308] ^ 11);
  assign w249[1] = |(datain[307:304] ^ 9);
  assign w249[2] = |(datain[303:300] ^ 11);
  assign w249[3] = |(datain[299:296] ^ 8);
  assign w249[4] = |(datain[295:292] ^ 0);
  assign w249[5] = |(datain[291:288] ^ 1);
  assign w249[6] = |(datain[287:284] ^ 8);
  assign w249[7] = |(datain[283:280] ^ 11);
  assign w249[8] = |(datain[279:276] ^ 13);
  assign w249[9] = |(datain[275:272] ^ 6);
  assign w249[10] = |(datain[271:268] ^ 12);
  assign w249[11] = |(datain[267:264] ^ 13);
  assign w249[12] = |(datain[263:260] ^ 2);
  assign w249[13] = |(datain[259:256] ^ 1);
  assign w249[14] = |(datain[255:252] ^ 7);
  assign w249[15] = |(datain[251:248] ^ 2);
  assign w249[16] = |(datain[247:244] ^ 1);
  assign w249[17] = |(datain[243:240] ^ 15);
  assign w249[18] = |(datain[239:236] ^ 3);
  assign w249[19] = |(datain[235:232] ^ 3);
  assign w249[20] = |(datain[231:228] ^ 13);
  assign w249[21] = |(datain[227:224] ^ 2);
  assign w249[22] = |(datain[223:220] ^ 3);
  assign w249[23] = |(datain[219:216] ^ 3);
  assign w249[24] = |(datain[215:212] ^ 12);
  assign w249[25] = |(datain[211:208] ^ 9);
  assign w249[26] = |(datain[207:204] ^ 11);
  assign w249[27] = |(datain[203:200] ^ 8);
  assign w249[28] = |(datain[199:196] ^ 0);
  assign w249[29] = |(datain[195:192] ^ 0);
  assign w249[30] = |(datain[191:188] ^ 4);
  assign w249[31] = |(datain[187:184] ^ 2);
  assign w249[32] = |(datain[183:180] ^ 12);
  assign w249[33] = |(datain[179:176] ^ 13);
  assign w249[34] = |(datain[175:172] ^ 2);
  assign w249[35] = |(datain[171:168] ^ 1);
  assign w249[36] = |(datain[167:164] ^ 7);
  assign w249[37] = |(datain[163:160] ^ 2);
  assign w249[38] = |(datain[159:156] ^ 1);
  assign w249[39] = |(datain[155:152] ^ 4);
  assign w249[40] = |(datain[151:148] ^ 2);
  assign w249[41] = |(datain[147:144] ^ 14);
  assign w249[42] = |(datain[143:140] ^ 10);
  assign w249[43] = |(datain[139:136] ^ 1);
  assign w249[44] = |(datain[135:132] ^ 9);
  assign w249[45] = |(datain[131:128] ^ 10);
  assign w249[46] = |(datain[127:124] ^ 0);
  assign w249[47] = |(datain[123:120] ^ 0);
  assign w249[48] = |(datain[119:116] ^ 12);
  assign w249[49] = |(datain[115:112] ^ 7);
  assign w249[50] = |(datain[111:108] ^ 0);
  assign w249[51] = |(datain[107:104] ^ 5);
  assign w249[52] = |(datain[103:100] ^ 4);
  assign w249[53] = |(datain[99:96] ^ 13);
  assign w249[54] = |(datain[95:92] ^ 14);
  assign w249[55] = |(datain[91:88] ^ 9);
  assign w249[56] = |(datain[87:84] ^ 8);
  assign w249[57] = |(datain[83:80] ^ 9);
  assign w249[58] = |(datain[79:76] ^ 4);
  assign w249[59] = |(datain[75:72] ^ 5);
  assign w249[60] = |(datain[71:68] ^ 0);
  assign w249[61] = |(datain[67:64] ^ 2);
  assign w249[62] = |(datain[63:60] ^ 11);
  assign w249[63] = |(datain[59:56] ^ 4);
  assign w249[64] = |(datain[55:52] ^ 4);
  assign w249[65] = |(datain[51:48] ^ 0);
  assign w249[66] = |(datain[47:44] ^ 11);
  assign w249[67] = |(datain[43:40] ^ 9);
  assign w249[68] = |(datain[39:36] ^ 0);
  assign w249[69] = |(datain[35:32] ^ 4);
  assign w249[70] = |(datain[31:28] ^ 0);
  assign w249[71] = |(datain[27:24] ^ 0);
  assign w249[72] = |(datain[23:20] ^ 8);
  assign w249[73] = |(datain[19:16] ^ 11);
  assign w249[74] = |(datain[15:12] ^ 13);
  assign w249[75] = |(datain[11:8] ^ 7);
  assign comp[249] = ~(|w249);
  wire [30-1:0] w250;
  assign w250[0] = |(datain[311:308] ^ 8);
  assign w250[1] = |(datain[307:304] ^ 11);
  assign w250[2] = |(datain[303:300] ^ 0);
  assign w250[3] = |(datain[299:296] ^ 1);
  assign w250[4] = |(datain[295:292] ^ 0);
  assign w250[5] = |(datain[291:288] ^ 3);
  assign w250[6] = |(datain[287:284] ^ 15);
  assign w250[7] = |(datain[283:280] ^ 5);
  assign w250[8] = |(datain[279:276] ^ 11);
  assign w250[9] = |(datain[275:272] ^ 15);
  assign w250[10] = |(datain[271:268] ^ 0);
  assign w250[11] = |(datain[267:264] ^ 0);
  assign w250[12] = |(datain[263:260] ^ 0);
  assign w250[13] = |(datain[259:256] ^ 1);
  assign w250[14] = |(datain[255:252] ^ 10);
  assign w250[15] = |(datain[251:248] ^ 5);
  assign w250[16] = |(datain[247:244] ^ 10);
  assign w250[17] = |(datain[243:240] ^ 5);
  assign w250[18] = |(datain[239:236] ^ 11);
  assign w250[19] = |(datain[235:232] ^ 8);
  assign w250[20] = |(datain[231:228] ^ 0);
  assign w250[21] = |(datain[227:224] ^ 0);
  assign w250[22] = |(datain[223:220] ^ 3);
  assign w250[23] = |(datain[219:216] ^ 3);
  assign w250[24] = |(datain[215:212] ^ 12);
  assign w250[25] = |(datain[211:208] ^ 13);
  assign w250[26] = |(datain[207:204] ^ 2);
  assign w250[27] = |(datain[203:200] ^ 1);
  assign w250[28] = |(datain[199:196] ^ 5);
  assign w250[29] = |(datain[195:192] ^ 2);
  assign comp[250] = ~(|w250);
  wire [46-1:0] w251;
  assign w251[0] = |(datain[311:308] ^ 12);
  assign w251[1] = |(datain[307:304] ^ 13);
  assign w251[2] = |(datain[303:300] ^ 2);
  assign w251[3] = |(datain[299:296] ^ 1);
  assign w251[4] = |(datain[295:292] ^ 11);
  assign w251[5] = |(datain[291:288] ^ 8);
  assign w251[6] = |(datain[287:284] ^ 2);
  assign w251[7] = |(datain[283:280] ^ 4);
  assign w251[8] = |(datain[279:276] ^ 3);
  assign w251[9] = |(datain[275:272] ^ 5);
  assign w251[10] = |(datain[271:268] ^ 12);
  assign w251[11] = |(datain[267:264] ^ 13);
  assign w251[12] = |(datain[263:260] ^ 2);
  assign w251[13] = |(datain[259:256] ^ 1);
  assign w251[14] = |(datain[255:252] ^ 5);
  assign w251[15] = |(datain[251:248] ^ 3);
  assign w251[16] = |(datain[247:244] ^ 0);
  assign w251[17] = |(datain[243:240] ^ 6);
  assign w251[18] = |(datain[239:236] ^ 11);
  assign w251[19] = |(datain[235:232] ^ 10);
  assign w251[20] = |(datain[231:228] ^ 1);
  assign w251[21] = |(datain[227:224] ^ 3);
  assign w251[22] = |(datain[223:220] ^ 0);
  assign w251[23] = |(datain[219:216] ^ 2);
  assign w251[24] = |(datain[215:212] ^ 0);
  assign w251[25] = |(datain[211:208] ^ 3);
  assign w251[26] = |(datain[207:204] ^ 13);
  assign w251[27] = |(datain[203:200] ^ 5);
  assign w251[28] = |(datain[199:196] ^ 11);
  assign w251[29] = |(datain[195:192] ^ 8);
  assign w251[30] = |(datain[191:188] ^ 2);
  assign w251[31] = |(datain[187:184] ^ 4);
  assign w251[32] = |(datain[183:180] ^ 2);
  assign w251[33] = |(datain[179:176] ^ 5);
  assign w251[34] = |(datain[175:172] ^ 12);
  assign w251[35] = |(datain[171:168] ^ 13);
  assign w251[36] = |(datain[167:164] ^ 2);
  assign w251[37] = |(datain[163:160] ^ 1);
  assign w251[38] = |(datain[159:156] ^ 8);
  assign w251[39] = |(datain[155:152] ^ 13);
  assign w251[40] = |(datain[151:148] ^ 9);
  assign w251[41] = |(datain[147:144] ^ 6);
  assign w251[42] = |(datain[143:140] ^ 5);
  assign w251[43] = |(datain[139:136] ^ 0);
  assign w251[44] = |(datain[135:132] ^ 0);
  assign w251[45] = |(datain[131:128] ^ 2);
  assign comp[251] = ~(|w251);
  wire [26-1:0] w252;
  assign w252[0] = |(datain[311:308] ^ 5);
  assign w252[1] = |(datain[307:304] ^ 1);
  assign w252[2] = |(datain[303:300] ^ 10);
  assign w252[3] = |(datain[299:296] ^ 13);
  assign w252[4] = |(datain[295:292] ^ 3);
  assign w252[5] = |(datain[291:288] ^ 3);
  assign w252[6] = |(datain[287:284] ^ 13);
  assign w252[7] = |(datain[283:280] ^ 0);
  assign w252[8] = |(datain[279:276] ^ 14);
  assign w252[9] = |(datain[275:272] ^ 2);
  assign w252[10] = |(datain[271:268] ^ 15);
  assign w252[11] = |(datain[267:264] ^ 11);
  assign w252[12] = |(datain[263:260] ^ 5);
  assign w252[13] = |(datain[259:256] ^ 9);
  assign w252[14] = |(datain[255:252] ^ 3);
  assign w252[15] = |(datain[251:248] ^ 1);
  assign w252[16] = |(datain[247:244] ^ 1);
  assign w252[17] = |(datain[243:240] ^ 5);
  assign w252[18] = |(datain[239:236] ^ 4);
  assign w252[19] = |(datain[235:232] ^ 7);
  assign w252[20] = |(datain[231:228] ^ 4);
  assign w252[21] = |(datain[227:224] ^ 7);
  assign w252[22] = |(datain[223:220] ^ 14);
  assign w252[23] = |(datain[219:216] ^ 2);
  assign w252[24] = |(datain[215:212] ^ 15);
  assign w252[25] = |(datain[211:208] ^ 10);
  assign comp[252] = ~(|w252);
  wire [32-1:0] w253;
  assign w253[0] = |(datain[311:308] ^ 11);
  assign w253[1] = |(datain[307:304] ^ 9);
  assign w253[2] = |(datain[303:300] ^ 8);
  assign w253[3] = |(datain[299:296] ^ 1);
  assign w253[4] = |(datain[295:292] ^ 0);
  assign w253[5] = |(datain[291:288] ^ 1);
  assign w253[6] = |(datain[287:284] ^ 5);
  assign w253[7] = |(datain[283:280] ^ 1);
  assign w253[8] = |(datain[279:276] ^ 10);
  assign w253[9] = |(datain[275:272] ^ 13);
  assign w253[10] = |(datain[271:268] ^ 3);
  assign w253[11] = |(datain[267:264] ^ 3);
  assign w253[12] = |(datain[263:260] ^ 13);
  assign w253[13] = |(datain[259:256] ^ 0);
  assign w253[14] = |(datain[255:252] ^ 14);
  assign w253[15] = |(datain[251:248] ^ 2);
  assign w253[16] = |(datain[247:244] ^ 15);
  assign w253[17] = |(datain[243:240] ^ 11);
  assign w253[18] = |(datain[239:236] ^ 5);
  assign w253[19] = |(datain[235:232] ^ 9);
  assign w253[20] = |(datain[231:228] ^ 3);
  assign w253[21] = |(datain[227:224] ^ 1);
  assign w253[22] = |(datain[223:220] ^ 1);
  assign w253[23] = |(datain[219:216] ^ 5);
  assign w253[24] = |(datain[215:212] ^ 4);
  assign w253[25] = |(datain[211:208] ^ 7);
  assign w253[26] = |(datain[207:204] ^ 4);
  assign w253[27] = |(datain[203:200] ^ 7);
  assign w253[28] = |(datain[199:196] ^ 14);
  assign w253[29] = |(datain[195:192] ^ 2);
  assign w253[30] = |(datain[191:188] ^ 15);
  assign w253[31] = |(datain[187:184] ^ 10);
  assign comp[253] = ~(|w253);
  wire [28-1:0] w254;
  assign w254[0] = |(datain[311:308] ^ 0);
  assign w254[1] = |(datain[307:304] ^ 6);
  assign w254[2] = |(datain[303:300] ^ 13);
  assign w254[3] = |(datain[299:296] ^ 4);
  assign w254[4] = |(datain[295:292] ^ 0);
  assign w254[5] = |(datain[291:288] ^ 3);
  assign w254[6] = |(datain[287:284] ^ 0);
  assign w254[7] = |(datain[283:280] ^ 1);
  assign w254[8] = |(datain[279:276] ^ 7);
  assign w254[9] = |(datain[275:272] ^ 4);
  assign w254[10] = |(datain[271:268] ^ 0);
  assign w254[11] = |(datain[267:264] ^ 7);
  assign w254[12] = |(datain[263:260] ^ 8);
  assign w254[13] = |(datain[259:256] ^ 14);
  assign w254[14] = |(datain[255:252] ^ 13);
  assign w254[15] = |(datain[251:248] ^ 0);
  assign w254[16] = |(datain[247:244] ^ 5);
  assign w254[17] = |(datain[243:240] ^ 3);
  assign w254[18] = |(datain[239:236] ^ 1);
  assign w254[19] = |(datain[235:232] ^ 14);
  assign w254[20] = |(datain[231:228] ^ 1);
  assign w254[21] = |(datain[227:224] ^ 14);
  assign w254[22] = |(datain[223:220] ^ 14);
  assign w254[23] = |(datain[219:216] ^ 11);
  assign w254[24] = |(datain[215:212] ^ 0);
  assign w254[25] = |(datain[211:208] ^ 5);
  assign w254[26] = |(datain[207:204] ^ 5);
  assign w254[27] = |(datain[203:200] ^ 0);
  assign comp[254] = ~(|w254);
  wire [32-1:0] w255;
  assign w255[0] = |(datain[311:308] ^ 1);
  assign w255[1] = |(datain[307:304] ^ 14);
  assign w255[2] = |(datain[303:300] ^ 6);
  assign w255[3] = |(datain[299:296] ^ 12);
  assign w255[4] = |(datain[295:292] ^ 0);
  assign w255[5] = |(datain[291:288] ^ 4);
  assign w255[6] = |(datain[287:284] ^ 8);
  assign w255[7] = |(datain[283:280] ^ 9);
  assign w255[8] = |(datain[279:276] ^ 1);
  assign w255[9] = |(datain[275:272] ^ 14);
  assign w255[10] = |(datain[271:268] ^ 6);
  assign w255[11] = |(datain[267:264] ^ 6);
  assign w255[12] = |(datain[263:260] ^ 0);
  assign w255[13] = |(datain[259:256] ^ 4);
  assign w255[14] = |(datain[255:252] ^ 0);
  assign w255[15] = |(datain[251:248] ^ 7);
  assign w255[16] = |(datain[247:244] ^ 11);
  assign w255[17] = |(datain[243:240] ^ 4);
  assign w255[18] = |(datain[239:236] ^ 1);
  assign w255[19] = |(datain[235:232] ^ 10);
  assign w255[20] = |(datain[231:228] ^ 11);
  assign w255[21] = |(datain[227:224] ^ 10);
  assign w255[22] = |(datain[223:220] ^ 6);
  assign w255[23] = |(datain[219:216] ^ 12);
  assign w255[24] = |(datain[215:212] ^ 0);
  assign w255[25] = |(datain[211:208] ^ 4);
  assign w255[26] = |(datain[207:204] ^ 12);
  assign w255[27] = |(datain[203:200] ^ 13);
  assign w255[28] = |(datain[199:196] ^ 2);
  assign w255[29] = |(datain[195:192] ^ 1);
  assign w255[30] = |(datain[191:188] ^ 12);
  assign w255[31] = |(datain[187:184] ^ 7);
  assign comp[255] = ~(|w255);
  wire [30-1:0] w256;
  assign w256[0] = |(datain[311:308] ^ 0);
  assign w256[1] = |(datain[307:304] ^ 4);
  assign w256[2] = |(datain[303:300] ^ 8);
  assign w256[3] = |(datain[299:296] ^ 1);
  assign w256[4] = |(datain[295:292] ^ 14);
  assign w256[5] = |(datain[291:288] ^ 1);
  assign w256[6] = |(datain[287:284] ^ 15);
  assign w256[7] = |(datain[283:280] ^ 8);
  assign w256[8] = |(datain[279:276] ^ 0);
  assign w256[9] = |(datain[275:272] ^ 0);
  assign w256[10] = |(datain[271:268] ^ 14);
  assign w256[11] = |(datain[267:264] ^ 8);
  assign w256[12] = |(datain[263:260] ^ 13);
  assign w256[13] = |(datain[259:256] ^ 1);
  assign w256[14] = |(datain[255:252] ^ 0);
  assign w256[15] = |(datain[251:248] ^ 1);
  assign w256[16] = |(datain[247:244] ^ 11);
  assign w256[17] = |(datain[243:240] ^ 8);
  assign w256[18] = |(datain[239:236] ^ 0);
  assign w256[19] = |(datain[235:232] ^ 2);
  assign w256[20] = |(datain[231:228] ^ 3);
  assign w256[21] = |(datain[227:224] ^ 13);
  assign w256[22] = |(datain[223:220] ^ 11);
  assign w256[23] = |(datain[219:216] ^ 10);
  assign w256[24] = |(datain[215:212] ^ 9);
  assign w256[25] = |(datain[211:208] ^ 6);
  assign w256[26] = |(datain[207:204] ^ 0);
  assign w256[27] = |(datain[203:200] ^ 4);
  assign w256[28] = |(datain[199:196] ^ 12);
  assign w256[29] = |(datain[195:192] ^ 13);
  assign comp[256] = ~(|w256);
  wire [42-1:0] w257;
  assign w257[0] = |(datain[311:308] ^ 4);
  assign w257[1] = |(datain[307:304] ^ 9);
  assign w257[2] = |(datain[303:300] ^ 11);
  assign w257[3] = |(datain[299:296] ^ 7);
  assign w257[4] = |(datain[295:292] ^ 4);
  assign w257[5] = |(datain[291:288] ^ 2);
  assign w257[6] = |(datain[287:284] ^ 4);
  assign w257[7] = |(datain[283:280] ^ 7);
  assign w257[8] = |(datain[279:276] ^ 3);
  assign w257[9] = |(datain[275:272] ^ 10);
  assign w257[10] = |(datain[271:268] ^ 2);
  assign w257[11] = |(datain[267:264] ^ 5);
  assign w257[12] = |(datain[263:260] ^ 7);
  assign w257[13] = |(datain[259:256] ^ 5);
  assign w257[14] = |(datain[255:252] ^ 1);
  assign w257[15] = |(datain[251:248] ^ 5);
  assign w257[16] = |(datain[247:244] ^ 3);
  assign w257[17] = |(datain[243:240] ^ 10);
  assign w257[18] = |(datain[239:236] ^ 7);
  assign w257[19] = |(datain[235:232] ^ 13);
  assign w257[20] = |(datain[231:228] ^ 0);
  assign w257[21] = |(datain[227:224] ^ 1);
  assign w257[22] = |(datain[223:220] ^ 7);
  assign w257[23] = |(datain[219:216] ^ 5);
  assign w257[24] = |(datain[215:212] ^ 1);
  assign w257[25] = |(datain[211:208] ^ 0);
  assign w257[26] = |(datain[207:204] ^ 3);
  assign w257[27] = |(datain[203:200] ^ 10);
  assign w257[28] = |(datain[199:196] ^ 4);
  assign w257[29] = |(datain[195:192] ^ 5);
  assign w257[30] = |(datain[191:188] ^ 0);
  assign w257[31] = |(datain[187:184] ^ 2);
  assign w257[32] = |(datain[183:180] ^ 7);
  assign w257[33] = |(datain[179:176] ^ 5);
  assign w257[34] = |(datain[175:172] ^ 0);
  assign w257[35] = |(datain[171:168] ^ 11);
  assign w257[36] = |(datain[167:164] ^ 12);
  assign w257[37] = |(datain[163:160] ^ 6);
  assign w257[38] = |(datain[159:156] ^ 4);
  assign w257[39] = |(datain[155:152] ^ 5);
  assign w257[40] = |(datain[151:148] ^ 0);
  assign w257[41] = |(datain[147:144] ^ 2);
  assign comp[257] = ~(|w257);
  wire [46-1:0] w258;
  assign w258[0] = |(datain[311:308] ^ 1);
  assign w258[1] = |(datain[307:304] ^ 1);
  assign w258[2] = |(datain[303:300] ^ 5);
  assign w258[3] = |(datain[299:296] ^ 11);
  assign w258[4] = |(datain[295:292] ^ 5);
  assign w258[5] = |(datain[291:288] ^ 9);
  assign w258[6] = |(datain[287:284] ^ 5);
  assign w258[7] = |(datain[283:280] ^ 10);
  assign w258[8] = |(datain[279:276] ^ 14);
  assign w258[9] = |(datain[275:272] ^ 8);
  assign w258[10] = |(datain[271:268] ^ 0);
  assign w258[11] = |(datain[267:264] ^ 0);
  assign w258[12] = |(datain[263:260] ^ 0);
  assign w258[13] = |(datain[259:256] ^ 0);
  assign w258[14] = |(datain[255:252] ^ 5);
  assign w258[15] = |(datain[251:248] ^ 13);
  assign w258[16] = |(datain[247:244] ^ 8);
  assign w258[17] = |(datain[243:240] ^ 1);
  assign w258[18] = |(datain[239:236] ^ 14);
  assign w258[19] = |(datain[235:232] ^ 13);
  assign w258[20] = |(datain[231:228] ^ 0);
  assign w258[21] = |(datain[227:224] ^ 11);
  assign w258[22] = |(datain[223:220] ^ 0);
  assign w258[23] = |(datain[219:216] ^ 0);
  assign w258[24] = |(datain[215:212] ^ 11);
  assign w258[25] = |(datain[211:208] ^ 8);
  assign w258[26] = |(datain[207:204] ^ 7);
  assign w258[27] = |(datain[203:200] ^ 7);
  assign w258[28] = |(datain[199:196] ^ 7);
  assign w258[29] = |(datain[195:192] ^ 7);
  assign w258[30] = |(datain[191:188] ^ 12);
  assign w258[31] = |(datain[187:184] ^ 13);
  assign w258[32] = |(datain[183:180] ^ 2);
  assign w258[33] = |(datain[179:176] ^ 1);
  assign w258[34] = |(datain[175:172] ^ 3);
  assign w258[35] = |(datain[171:168] ^ 13);
  assign w258[36] = |(datain[167:164] ^ 8);
  assign w258[37] = |(datain[163:160] ^ 8);
  assign w258[38] = |(datain[159:156] ^ 8);
  assign w258[39] = |(datain[155:152] ^ 8);
  assign w258[40] = |(datain[151:148] ^ 7);
  assign w258[41] = |(datain[147:144] ^ 4);
  assign w258[42] = |(datain[143:140] ^ 5);
  assign w258[43] = |(datain[139:136] ^ 12);
  assign w258[44] = |(datain[135:132] ^ 11);
  assign w258[45] = |(datain[131:128] ^ 4);
  assign comp[258] = ~(|w258);
  wire [36-1:0] w259;
  assign w259[0] = |(datain[311:308] ^ 4);
  assign w259[1] = |(datain[307:304] ^ 4);
  assign w259[2] = |(datain[303:300] ^ 5);
  assign w259[3] = |(datain[299:296] ^ 11);
  assign w259[4] = |(datain[295:292] ^ 7);
  assign w259[5] = |(datain[291:288] ^ 2);
  assign w259[6] = |(datain[287:284] ^ 1);
  assign w259[7] = |(datain[283:280] ^ 9);
  assign w259[8] = |(datain[279:276] ^ 11);
  assign w259[9] = |(datain[275:272] ^ 8);
  assign w259[10] = |(datain[271:268] ^ 9);
  assign w259[11] = |(datain[267:264] ^ 0);
  assign w259[12] = |(datain[263:260] ^ 7);
  assign w259[13] = |(datain[259:256] ^ 14);
  assign w259[14] = |(datain[255:252] ^ 14);
  assign w259[15] = |(datain[251:248] ^ 8);
  assign w259[16] = |(datain[247:244] ^ 12);
  assign w259[17] = |(datain[243:240] ^ 8);
  assign w259[18] = |(datain[239:236] ^ 0);
  assign w259[19] = |(datain[235:232] ^ 0);
  assign w259[20] = |(datain[231:228] ^ 11);
  assign w259[21] = |(datain[227:224] ^ 8);
  assign w259[22] = |(datain[223:220] ^ 0);
  assign w259[23] = |(datain[219:216] ^ 8);
  assign w259[24] = |(datain[215:212] ^ 3);
  assign w259[25] = |(datain[211:208] ^ 5);
  assign w259[26] = |(datain[207:204] ^ 12);
  assign w259[27] = |(datain[203:200] ^ 13);
  assign w259[28] = |(datain[199:196] ^ 2);
  assign w259[29] = |(datain[195:192] ^ 1);
  assign w259[30] = |(datain[191:188] ^ 8);
  assign w259[31] = |(datain[187:184] ^ 9);
  assign w259[32] = |(datain[183:180] ^ 5);
  assign w259[33] = |(datain[179:176] ^ 12);
  assign w259[34] = |(datain[175:172] ^ 5);
  assign w259[35] = |(datain[171:168] ^ 13);
  assign comp[259] = ~(|w259);
  wire [32-1:0] w260;
  assign w260[0] = |(datain[311:308] ^ 0);
  assign w260[1] = |(datain[307:304] ^ 15);
  assign w260[2] = |(datain[303:300] ^ 14);
  assign w260[3] = |(datain[299:296] ^ 0);
  assign w260[4] = |(datain[295:292] ^ 12);
  assign w260[5] = |(datain[291:288] ^ 13);
  assign w260[6] = |(datain[287:284] ^ 2);
  assign w260[7] = |(datain[283:280] ^ 1);
  assign w260[8] = |(datain[279:276] ^ 3);
  assign w260[9] = |(datain[275:272] ^ 13);
  assign w260[10] = |(datain[271:268] ^ 3);
  assign w260[11] = |(datain[267:264] ^ 1);
  assign w260[12] = |(datain[263:260] ^ 4);
  assign w260[13] = |(datain[259:256] ^ 12);
  assign w260[14] = |(datain[255:252] ^ 7);
  assign w260[15] = |(datain[251:248] ^ 5);
  assign w260[16] = |(datain[247:244] ^ 3);
  assign w260[17] = |(datain[243:240] ^ 13);
  assign w260[18] = |(datain[239:236] ^ 2);
  assign w260[19] = |(datain[235:232] ^ 14);
  assign w260[20] = |(datain[231:228] ^ 8);
  assign w260[21] = |(datain[227:224] ^ 1);
  assign w260[22] = |(datain[223:220] ^ 3);
  assign w260[23] = |(datain[219:216] ^ 14);
  assign w260[24] = |(datain[215:212] ^ 2);
  assign w260[25] = |(datain[211:208] ^ 11);
  assign w260[26] = |(datain[207:204] ^ 0);
  assign w260[27] = |(datain[203:200] ^ 0);
  assign w260[28] = |(datain[199:196] ^ 4);
  assign w260[29] = |(datain[195:192] ^ 13);
  assign w260[30] = |(datain[191:188] ^ 5);
  assign w260[31] = |(datain[187:184] ^ 10);
  assign comp[260] = ~(|w260);
  wire [30-1:0] w261;
  assign w261[0] = |(datain[311:308] ^ 8);
  assign w261[1] = |(datain[307:304] ^ 14);
  assign w261[2] = |(datain[303:300] ^ 12);
  assign w261[3] = |(datain[299:296] ^ 0);
  assign w261[4] = |(datain[295:292] ^ 8);
  assign w261[5] = |(datain[291:288] ^ 14);
  assign w261[6] = |(datain[287:284] ^ 13);
  assign w261[7] = |(datain[283:280] ^ 8);
  assign w261[8] = |(datain[279:276] ^ 8);
  assign w261[9] = |(datain[275:272] ^ 0);
  assign w261[10] = |(datain[271:268] ^ 3);
  assign w261[11] = |(datain[267:264] ^ 14);
  assign w261[12] = |(datain[263:260] ^ 0);
  assign w261[13] = |(datain[259:256] ^ 0);
  assign w261[14] = |(datain[255:252] ^ 0);
  assign w261[15] = |(datain[251:248] ^ 0);
  assign w261[16] = |(datain[247:244] ^ 5);
  assign w261[17] = |(datain[243:240] ^ 10);
  assign w261[18] = |(datain[239:236] ^ 7);
  assign w261[19] = |(datain[235:232] ^ 4);
  assign w261[20] = |(datain[231:228] ^ 1);
  assign w261[21] = |(datain[227:224] ^ 5);
  assign w261[22] = |(datain[223:220] ^ 0);
  assign w261[23] = |(datain[219:216] ^ 3);
  assign w261[24] = |(datain[215:212] ^ 0);
  assign w261[25] = |(datain[211:208] ^ 6);
  assign w261[26] = |(datain[207:204] ^ 0);
  assign w261[27] = |(datain[203:200] ^ 3);
  assign w261[28] = |(datain[199:196] ^ 0);
  assign w261[29] = |(datain[195:192] ^ 0);
  assign comp[261] = ~(|w261);
  wire [44-1:0] w262;
  assign w262[0] = |(datain[311:308] ^ 0);
  assign w262[1] = |(datain[307:304] ^ 3);
  assign w262[2] = |(datain[303:300] ^ 5);
  assign w262[3] = |(datain[299:296] ^ 3);
  assign w262[4] = |(datain[295:292] ^ 2);
  assign w262[5] = |(datain[291:288] ^ 14);
  assign w262[6] = |(datain[287:284] ^ 15);
  assign w262[7] = |(datain[283:280] ^ 15);
  assign w262[8] = |(datain[279:276] ^ 11);
  assign w262[9] = |(datain[275:272] ^ 5);
  assign w262[10] = |(datain[271:268] ^ 5);
  assign w262[11] = |(datain[267:264] ^ 13);
  assign w262[12] = |(datain[263:260] ^ 0);
  assign w262[13] = |(datain[259:256] ^ 4);
  assign w262[14] = |(datain[255:252] ^ 11);
  assign w262[15] = |(datain[251:248] ^ 11);
  assign w262[16] = |(datain[247:244] ^ 13);
  assign w262[17] = |(datain[243:240] ^ 14);
  assign w262[18] = |(datain[239:236] ^ 0);
  assign w262[19] = |(datain[235:232] ^ 3);
  assign w262[20] = |(datain[231:228] ^ 11);
  assign w262[21] = |(datain[227:224] ^ 9);
  assign w262[22] = |(datain[223:220] ^ 7);
  assign w262[23] = |(datain[219:216] ^ 15);
  assign w262[24] = |(datain[215:212] ^ 0);
  assign w262[25] = |(datain[211:208] ^ 0);
  assign w262[26] = |(datain[207:204] ^ 5);
  assign w262[27] = |(datain[203:200] ^ 8);
  assign w262[28] = |(datain[199:196] ^ 2);
  assign w262[29] = |(datain[195:192] ^ 14);
  assign w262[30] = |(datain[191:188] ^ 3);
  assign w262[31] = |(datain[187:184] ^ 0);
  assign w262[32] = |(datain[183:180] ^ 0);
  assign w262[33] = |(datain[179:176] ^ 1);
  assign w262[34] = |(datain[175:172] ^ 4);
  assign w262[35] = |(datain[171:168] ^ 3);
  assign w262[36] = |(datain[167:164] ^ 14);
  assign w262[37] = |(datain[163:160] ^ 2);
  assign w262[38] = |(datain[159:156] ^ 15);
  assign w262[39] = |(datain[155:152] ^ 10);
  assign w262[40] = |(datain[151:148] ^ 5);
  assign w262[41] = |(datain[147:144] ^ 11);
  assign w262[42] = |(datain[143:140] ^ 14);
  assign w262[43] = |(datain[139:136] ^ 8);
  assign comp[262] = ~(|w262);
  wire [30-1:0] w263;
  assign w263[0] = |(datain[311:308] ^ 12);
  assign w263[1] = |(datain[307:304] ^ 7);
  assign w263[2] = |(datain[303:300] ^ 0);
  assign w263[3] = |(datain[299:296] ^ 3);
  assign w263[4] = |(datain[295:292] ^ 5);
  assign w263[5] = |(datain[291:288] ^ 3);
  assign w263[6] = |(datain[287:284] ^ 2);
  assign w263[7] = |(datain[283:280] ^ 14);
  assign w263[8] = |(datain[279:276] ^ 15);
  assign w263[9] = |(datain[275:272] ^ 15);
  assign w263[10] = |(datain[271:268] ^ 11);
  assign w263[11] = |(datain[267:264] ^ 5);
  assign w263[12] = |(datain[263:260] ^ 5);
  assign w263[13] = |(datain[259:256] ^ 13);
  assign w263[14] = |(datain[255:252] ^ 0);
  assign w263[15] = |(datain[251:248] ^ 4);
  assign w263[16] = |(datain[247:244] ^ 11);
  assign w263[17] = |(datain[243:240] ^ 11);
  assign w263[18] = |(datain[239:236] ^ 13);
  assign w263[19] = |(datain[235:232] ^ 14);
  assign w263[20] = |(datain[231:228] ^ 0);
  assign w263[21] = |(datain[227:224] ^ 3);
  assign w263[22] = |(datain[223:220] ^ 11);
  assign w263[23] = |(datain[219:216] ^ 9);
  assign w263[24] = |(datain[215:212] ^ 7);
  assign w263[25] = |(datain[211:208] ^ 15);
  assign w263[26] = |(datain[207:204] ^ 0);
  assign w263[27] = |(datain[203:200] ^ 0);
  assign w263[28] = |(datain[199:196] ^ 5);
  assign w263[29] = |(datain[195:192] ^ 8);
  assign comp[263] = ~(|w263);
  wire [36-1:0] w264;
  assign w264[0] = |(datain[311:308] ^ 0);
  assign w264[1] = |(datain[307:304] ^ 3);
  assign w264[2] = |(datain[303:300] ^ 0);
  assign w264[3] = |(datain[299:296] ^ 3);
  assign w264[4] = |(datain[295:292] ^ 11);
  assign w264[5] = |(datain[291:288] ^ 4);
  assign w264[6] = |(datain[287:284] ^ 4);
  assign w264[7] = |(datain[283:280] ^ 0);
  assign w264[8] = |(datain[279:276] ^ 11);
  assign w264[9] = |(datain[275:272] ^ 9);
  assign w264[10] = |(datain[271:268] ^ 0);
  assign w264[11] = |(datain[267:264] ^ 3);
  assign w264[12] = |(datain[263:260] ^ 0);
  assign w264[13] = |(datain[259:256] ^ 0);
  assign w264[14] = |(datain[255:252] ^ 11);
  assign w264[15] = |(datain[251:248] ^ 10);
  assign w264[16] = |(datain[247:244] ^ 1);
  assign w264[17] = |(datain[243:240] ^ 6);
  assign w264[18] = |(datain[239:236] ^ 0);
  assign w264[19] = |(datain[235:232] ^ 3);
  assign w264[20] = |(datain[231:228] ^ 12);
  assign w264[21] = |(datain[227:224] ^ 13);
  assign w264[22] = |(datain[223:220] ^ 2);
  assign w264[23] = |(datain[219:216] ^ 1);
  assign w264[24] = |(datain[215:212] ^ 12);
  assign w264[25] = |(datain[211:208] ^ 3);
  assign w264[26] = |(datain[207:204] ^ 8);
  assign w264[27] = |(datain[203:200] ^ 11);
  assign w264[28] = |(datain[199:196] ^ 1);
  assign w264[29] = |(datain[195:192] ^ 14);
  assign w264[30] = |(datain[191:188] ^ 0);
  assign w264[31] = |(datain[187:184] ^ 8);
  assign w264[32] = |(datain[183:180] ^ 0);
  assign w264[33] = |(datain[179:176] ^ 3);
  assign w264[34] = |(datain[175:172] ^ 11);
  assign w264[35] = |(datain[171:168] ^ 8);
  assign comp[264] = ~(|w264);
  wire [32-1:0] w265;
  assign w265[0] = |(datain[311:308] ^ 14);
  assign w265[1] = |(datain[307:304] ^ 9);
  assign w265[2] = |(datain[303:300] ^ 10);
  assign w265[3] = |(datain[299:296] ^ 13);
  assign w265[4] = |(datain[295:292] ^ 0);
  assign w265[5] = |(datain[291:288] ^ 0);
  assign w265[6] = |(datain[287:284] ^ 11);
  assign w265[7] = |(datain[283:280] ^ 8);
  assign w265[8] = |(datain[279:276] ^ 11);
  assign w265[9] = |(datain[275:272] ^ 11);
  assign w265[10] = |(datain[271:268] ^ 11);
  assign w265[11] = |(datain[267:264] ^ 11);
  assign w265[12] = |(datain[263:260] ^ 12);
  assign w265[13] = |(datain[259:256] ^ 13);
  assign w265[14] = |(datain[255:252] ^ 2);
  assign w265[15] = |(datain[251:248] ^ 1);
  assign w265[16] = |(datain[247:244] ^ 3);
  assign w265[17] = |(datain[243:240] ^ 13);
  assign w265[18] = |(datain[239:236] ^ 6);
  assign w265[19] = |(datain[235:232] ^ 9);
  assign w265[20] = |(datain[231:228] ^ 6);
  assign w265[21] = |(datain[227:224] ^ 9);
  assign w265[22] = |(datain[223:220] ^ 7);
  assign w265[23] = |(datain[219:216] ^ 4);
  assign w265[24] = |(datain[215:212] ^ 0);
  assign w265[25] = |(datain[211:208] ^ 3);
  assign w265[26] = |(datain[207:204] ^ 14);
  assign w265[27] = |(datain[203:200] ^ 8);
  assign w265[28] = |(datain[199:196] ^ 3);
  assign w265[29] = |(datain[195:192] ^ 5);
  assign w265[30] = |(datain[191:188] ^ 0);
  assign w265[31] = |(datain[187:184] ^ 0);
  assign comp[265] = ~(|w265);
  wire [32-1:0] w266;
  assign w266[0] = |(datain[311:308] ^ 14);
  assign w266[1] = |(datain[307:304] ^ 8);
  assign w266[2] = |(datain[303:300] ^ 15);
  assign w266[3] = |(datain[299:296] ^ 15);
  assign w266[4] = |(datain[295:292] ^ 0);
  assign w266[5] = |(datain[291:288] ^ 0);
  assign w266[6] = |(datain[287:284] ^ 11);
  assign w266[7] = |(datain[283:280] ^ 4);
  assign w266[8] = |(datain[279:276] ^ 3);
  assign w266[9] = |(datain[275:272] ^ 15);
  assign w266[10] = |(datain[271:268] ^ 11);
  assign w266[11] = |(datain[267:264] ^ 9);
  assign w266[12] = |(datain[263:260] ^ 11);
  assign w266[13] = |(datain[259:256] ^ 9);
  assign w266[14] = |(datain[255:252] ^ 0);
  assign w266[15] = |(datain[251:248] ^ 3);
  assign w266[16] = |(datain[247:244] ^ 11);
  assign w266[17] = |(datain[243:240] ^ 10);
  assign w266[18] = |(datain[239:236] ^ 13);
  assign w266[19] = |(datain[235:232] ^ 5);
  assign w266[20] = |(datain[231:228] ^ 0);
  assign w266[21] = |(datain[227:224] ^ 4);
  assign w266[22] = |(datain[223:220] ^ 12);
  assign w266[23] = |(datain[219:216] ^ 13);
  assign w266[24] = |(datain[215:212] ^ 2);
  assign w266[25] = |(datain[211:208] ^ 1);
  assign w266[26] = |(datain[207:204] ^ 2);
  assign w266[27] = |(datain[203:200] ^ 10);
  assign w266[28] = |(datain[199:196] ^ 12);
  assign w266[29] = |(datain[195:192] ^ 0);
  assign w266[30] = |(datain[191:188] ^ 14);
  assign w266[31] = |(datain[187:184] ^ 8);
  assign comp[266] = ~(|w266);
  wire [46-1:0] w267;
  assign w267[0] = |(datain[311:308] ^ 6);
  assign w267[1] = |(datain[307:304] ^ 0);
  assign w267[2] = |(datain[303:300] ^ 3);
  assign w267[3] = |(datain[299:296] ^ 5);
  assign w267[4] = |(datain[295:292] ^ 12);
  assign w267[5] = |(datain[291:288] ^ 13);
  assign w267[6] = |(datain[287:284] ^ 2);
  assign w267[7] = |(datain[283:280] ^ 1);
  assign w267[8] = |(datain[279:276] ^ 8);
  assign w267[9] = |(datain[275:272] ^ 1);
  assign w267[10] = |(datain[271:268] ^ 15);
  assign w267[11] = |(datain[267:264] ^ 11);
  assign w267[12] = |(datain[263:260] ^ 3);
  assign w267[13] = |(datain[259:256] ^ 4);
  assign w267[14] = |(datain[255:252] ^ 1);
  assign w267[15] = |(datain[251:248] ^ 2);
  assign w267[16] = |(datain[247:244] ^ 7);
  assign w267[17] = |(datain[243:240] ^ 4);
  assign w267[18] = |(datain[239:236] ^ 0);
  assign w267[19] = |(datain[235:232] ^ 3);
  assign w267[20] = |(datain[231:228] ^ 14);
  assign w267[21] = |(datain[227:224] ^ 9);
  assign w267[22] = |(datain[223:220] ^ 12);
  assign w267[23] = |(datain[219:216] ^ 9);
  assign w267[24] = |(datain[215:212] ^ 0);
  assign w267[25] = |(datain[211:208] ^ 3);
  assign w267[26] = |(datain[207:204] ^ 14);
  assign w267[27] = |(datain[203:200] ^ 9);
  assign w267[28] = |(datain[199:196] ^ 0);
  assign w267[29] = |(datain[195:192] ^ 10);
  assign w267[30] = |(datain[191:188] ^ 0);
  assign w267[31] = |(datain[187:184] ^ 3);
  assign w267[32] = |(datain[183:180] ^ 5);
  assign w267[33] = |(datain[179:176] ^ 0);
  assign w267[34] = |(datain[175:172] ^ 5);
  assign w267[35] = |(datain[171:168] ^ 3);
  assign w267[36] = |(datain[167:164] ^ 5);
  assign w267[37] = |(datain[163:160] ^ 1);
  assign w267[38] = |(datain[159:156] ^ 5);
  assign w267[39] = |(datain[155:152] ^ 2);
  assign w267[40] = |(datain[151:148] ^ 1);
  assign w267[41] = |(datain[147:144] ^ 14);
  assign w267[42] = |(datain[143:140] ^ 0);
  assign w267[43] = |(datain[139:136] ^ 6);
  assign w267[44] = |(datain[135:132] ^ 5);
  assign w267[45] = |(datain[131:128] ^ 7);
  assign comp[267] = ~(|w267);
  wire [74-1:0] w268;
  assign w268[0] = |(datain[311:308] ^ 11);
  assign w268[1] = |(datain[307:304] ^ 8);
  assign w268[2] = |(datain[303:300] ^ 0);
  assign w268[3] = |(datain[299:296] ^ 12);
  assign w268[4] = |(datain[295:292] ^ 0);
  assign w268[5] = |(datain[291:288] ^ 2);
  assign w268[6] = |(datain[287:284] ^ 11);
  assign w268[7] = |(datain[283:280] ^ 9);
  assign w268[8] = |(datain[279:276] ^ 0);
  assign w268[9] = |(datain[275:272] ^ 3);
  assign w268[10] = |(datain[271:268] ^ 0);
  assign w268[11] = |(datain[267:264] ^ 0);
  assign w268[12] = |(datain[263:260] ^ 11);
  assign w268[13] = |(datain[259:256] ^ 10);
  assign w268[14] = |(datain[255:252] ^ 8);
  assign w268[15] = |(datain[251:248] ^ 0);
  assign w268[16] = |(datain[247:244] ^ 0);
  assign w268[17] = |(datain[243:240] ^ 0);
  assign w268[18] = |(datain[239:236] ^ 12);
  assign w268[19] = |(datain[235:232] ^ 13);
  assign w268[20] = |(datain[231:228] ^ 1);
  assign w268[21] = |(datain[227:224] ^ 3);
  assign w268[22] = |(datain[223:220] ^ 14);
  assign w268[23] = |(datain[219:216] ^ 11);
  assign w268[24] = |(datain[215:212] ^ 0);
  assign w268[25] = |(datain[211:208] ^ 2);
  assign w268[26] = |(datain[207:204] ^ 9);
  assign w268[27] = |(datain[203:200] ^ 0);
  assign w268[28] = |(datain[199:196] ^ 5);
  assign w268[29] = |(datain[195:192] ^ 6);
  assign w268[30] = |(datain[191:188] ^ 11);
  assign w268[31] = |(datain[187:184] ^ 4);
  assign w268[32] = |(datain[183:180] ^ 3);
  assign w268[33] = |(datain[179:176] ^ 0);
  assign w268[34] = |(datain[175:172] ^ 12);
  assign w268[35] = |(datain[171:168] ^ 13);
  assign w268[36] = |(datain[167:164] ^ 2);
  assign w268[37] = |(datain[163:160] ^ 1);
  assign w268[38] = |(datain[159:156] ^ 3);
  assign w268[39] = |(datain[155:152] ^ 12);
  assign w268[40] = |(datain[151:148] ^ 0);
  assign w268[41] = |(datain[147:144] ^ 3);
  assign w268[42] = |(datain[143:140] ^ 14);
  assign w268[43] = |(datain[139:136] ^ 11);
  assign w268[44] = |(datain[135:132] ^ 0);
  assign w268[45] = |(datain[131:128] ^ 1);
  assign w268[46] = |(datain[127:124] ^ 9);
  assign w268[47] = |(datain[123:120] ^ 0);
  assign w268[48] = |(datain[119:116] ^ 2);
  assign w268[49] = |(datain[115:112] ^ 14);
  assign w268[50] = |(datain[111:108] ^ 12);
  assign w268[51] = |(datain[107:104] ^ 6);
  assign w268[52] = |(datain[103:100] ^ 0);
  assign w268[53] = |(datain[99:96] ^ 6);
  assign w268[54] = |(datain[95:92] ^ 6);
  assign w268[55] = |(datain[91:88] ^ 2);
  assign w268[56] = |(datain[87:84] ^ 0);
  assign w268[57] = |(datain[83:80] ^ 2);
  assign w268[58] = |(datain[79:76] ^ 15);
  assign w268[59] = |(datain[75:72] ^ 15);
  assign w268[60] = |(datain[71:68] ^ 14);
  assign w268[61] = |(datain[67:64] ^ 8);
  assign w268[62] = |(datain[63:60] ^ 9);
  assign w268[63] = |(datain[59:56] ^ 0);
  assign w268[64] = |(datain[55:52] ^ 0);
  assign w268[65] = |(datain[51:48] ^ 2);
  assign w268[66] = |(datain[47:44] ^ 2);
  assign w268[67] = |(datain[43:40] ^ 14);
  assign w268[68] = |(datain[39:36] ^ 8);
  assign w268[69] = |(datain[35:32] ^ 0);
  assign w268[70] = |(datain[31:28] ^ 3);
  assign w268[71] = |(datain[27:24] ^ 14);
  assign w268[72] = |(datain[23:20] ^ 0);
  assign w268[73] = |(datain[19:16] ^ 15);
  assign comp[268] = ~(|w268);
  wire [76-1:0] w269;
  assign w269[0] = |(datain[311:308] ^ 11);
  assign w269[1] = |(datain[307:304] ^ 10);
  assign w269[2] = |(datain[303:300] ^ 0);
  assign w269[3] = |(datain[299:296] ^ 0);
  assign w269[4] = |(datain[295:292] ^ 0);
  assign w269[5] = |(datain[291:288] ^ 0);
  assign w269[6] = |(datain[287:284] ^ 11);
  assign w269[7] = |(datain[283:280] ^ 4);
  assign w269[8] = |(datain[279:276] ^ 4);
  assign w269[9] = |(datain[275:272] ^ 0);
  assign w269[10] = |(datain[271:268] ^ 12);
  assign w269[11] = |(datain[267:264] ^ 13);
  assign w269[12] = |(datain[263:260] ^ 2);
  assign w269[13] = |(datain[259:256] ^ 1);
  assign w269[14] = |(datain[255:252] ^ 14);
  assign w269[15] = |(datain[251:248] ^ 8);
  assign w269[16] = |(datain[247:244] ^ 7);
  assign w269[17] = |(datain[243:240] ^ 0);
  assign w269[18] = |(datain[239:236] ^ 0);
  assign w269[19] = |(datain[235:232] ^ 0);
  assign w269[20] = |(datain[231:228] ^ 11);
  assign w269[21] = |(datain[227:224] ^ 4);
  assign w269[22] = |(datain[223:220] ^ 3);
  assign w269[23] = |(datain[219:216] ^ 14);
  assign w269[24] = |(datain[215:212] ^ 12);
  assign w269[25] = |(datain[211:208] ^ 13);
  assign w269[26] = |(datain[207:204] ^ 2);
  assign w269[27] = |(datain[203:200] ^ 1);
  assign w269[28] = |(datain[199:196] ^ 12);
  assign w269[29] = |(datain[195:192] ^ 3);
  assign w269[30] = |(datain[191:188] ^ 11);
  assign w269[31] = |(datain[187:184] ^ 14);
  assign w269[32] = |(datain[183:180] ^ 0);
  assign w269[33] = |(datain[179:176] ^ 8);
  assign w269[34] = |(datain[175:172] ^ 0);
  assign w269[35] = |(datain[171:168] ^ 1);
  assign w269[36] = |(datain[167:164] ^ 11);
  assign w269[37] = |(datain[163:160] ^ 2);
  assign w269[38] = |(datain[159:156] ^ 0);
  assign w269[39] = |(datain[155:152] ^ 0);
  assign w269[40] = |(datain[151:148] ^ 11);
  assign w269[41] = |(datain[147:144] ^ 4);
  assign w269[42] = |(datain[143:140] ^ 4);
  assign w269[43] = |(datain[139:136] ^ 7);
  assign w269[44] = |(datain[135:132] ^ 12);
  assign w269[45] = |(datain[131:128] ^ 13);
  assign w269[46] = |(datain[127:124] ^ 2);
  assign w269[47] = |(datain[123:120] ^ 1);
  assign w269[48] = |(datain[119:116] ^ 12);
  assign w269[49] = |(datain[115:112] ^ 3);
  assign w269[50] = |(datain[111:108] ^ 0);
  assign w269[51] = |(datain[107:104] ^ 14);
  assign w269[52] = |(datain[103:100] ^ 1);
  assign w269[53] = |(datain[99:96] ^ 15);
  assign w269[54] = |(datain[95:92] ^ 11);
  assign w269[55] = |(datain[91:88] ^ 10);
  assign w269[56] = |(datain[87:84] ^ 4);
  assign w269[57] = |(datain[83:80] ^ 9);
  assign w269[58] = |(datain[79:76] ^ 0);
  assign w269[59] = |(datain[75:72] ^ 1);
  assign w269[60] = |(datain[71:68] ^ 11);
  assign w269[61] = |(datain[67:64] ^ 8);
  assign w269[62] = |(datain[63:60] ^ 0);
  assign w269[63] = |(datain[59:56] ^ 2);
  assign w269[64] = |(datain[55:52] ^ 3);
  assign w269[65] = |(datain[51:48] ^ 13);
  assign w269[66] = |(datain[47:44] ^ 12);
  assign w269[67] = |(datain[43:40] ^ 13);
  assign w269[68] = |(datain[39:36] ^ 2);
  assign w269[69] = |(datain[35:32] ^ 1);
  assign w269[70] = |(datain[31:28] ^ 5);
  assign w269[71] = |(datain[27:24] ^ 0);
  assign w269[72] = |(datain[23:20] ^ 5);
  assign w269[73] = |(datain[19:16] ^ 11);
  assign w269[74] = |(datain[15:12] ^ 12);
  assign w269[75] = |(datain[11:8] ^ 3);
  assign comp[269] = ~(|w269);
  wire [46-1:0] w270;
  assign w270[0] = |(datain[311:308] ^ 0);
  assign w270[1] = |(datain[307:304] ^ 5);
  assign w270[2] = |(datain[303:300] ^ 0);
  assign w270[3] = |(datain[299:296] ^ 5);
  assign w270[4] = |(datain[295:292] ^ 4);
  assign w270[5] = |(datain[291:288] ^ 7);
  assign w270[6] = |(datain[287:284] ^ 14);
  assign w270[7] = |(datain[283:280] ^ 2);
  assign w270[8] = |(datain[279:276] ^ 15);
  assign w270[9] = |(datain[275:272] ^ 10);
  assign w270[10] = |(datain[271:268] ^ 11);
  assign w270[11] = |(datain[267:264] ^ 9);
  assign w270[12] = |(datain[263:260] ^ 4);
  assign w270[13] = |(datain[259:256] ^ 12);
  assign w270[14] = |(datain[255:252] ^ 0);
  assign w270[15] = |(datain[251:248] ^ 4);
  assign w270[16] = |(datain[247:244] ^ 11);
  assign w270[17] = |(datain[243:240] ^ 10);
  assign w270[18] = |(datain[239:236] ^ 0);
  assign w270[19] = |(datain[235:232] ^ 0);
  assign w270[20] = |(datain[231:228] ^ 0);
  assign w270[21] = |(datain[227:224] ^ 0);
  assign w270[22] = |(datain[223:220] ^ 14);
  assign w270[23] = |(datain[219:216] ^ 8);
  assign w270[24] = |(datain[215:212] ^ 3);
  assign w270[25] = |(datain[211:208] ^ 8);
  assign w270[26] = |(datain[207:204] ^ 0);
  assign w270[27] = |(datain[203:200] ^ 0);
  assign w270[28] = |(datain[199:196] ^ 11);
  assign w270[29] = |(datain[195:192] ^ 15);
  assign w270[30] = |(datain[191:188] ^ 14);
  assign w270[31] = |(datain[187:184] ^ 11);
  assign w270[32] = |(datain[183:180] ^ 0);
  assign w270[33] = |(datain[179:176] ^ 1);
  assign w270[34] = |(datain[175:172] ^ 11);
  assign w270[35] = |(datain[171:168] ^ 9);
  assign w270[36] = |(datain[167:164] ^ 10);
  assign w270[37] = |(datain[163:160] ^ 0);
  assign w270[38] = |(datain[159:156] ^ 0);
  assign w270[39] = |(datain[155:152] ^ 0);
  assign w270[40] = |(datain[151:148] ^ 9);
  assign w270[41] = |(datain[147:144] ^ 12);
  assign w270[42] = |(datain[143:140] ^ 8);
  assign w270[43] = |(datain[139:136] ^ 0);
  assign w270[44] = |(datain[135:132] ^ 2);
  assign w270[45] = |(datain[131:128] ^ 13);
  assign comp[270] = ~(|w270);
  wire [42-1:0] w271;
  assign w271[0] = |(datain[311:308] ^ 8);
  assign w271[1] = |(datain[307:304] ^ 6);
  assign w271[2] = |(datain[303:300] ^ 0);
  assign w271[3] = |(datain[299:296] ^ 0);
  assign w271[4] = |(datain[295:292] ^ 8);
  assign w271[5] = |(datain[291:288] ^ 14);
  assign w271[6] = |(datain[287:284] ^ 12);
  assign w271[7] = |(datain[283:280] ^ 1);
  assign w271[8] = |(datain[279:276] ^ 2);
  assign w271[9] = |(datain[275:272] ^ 6);
  assign w271[10] = |(datain[271:268] ^ 8);
  assign w271[11] = |(datain[267:264] ^ 1);
  assign w271[12] = |(datain[263:260] ^ 7);
  assign w271[13] = |(datain[259:256] ^ 15);
  assign w271[14] = |(datain[255:252] ^ 0);
  assign w271[15] = |(datain[251:248] ^ 3);
  assign w271[16] = |(datain[247:244] ^ 4);
  assign w271[17] = |(datain[243:240] ^ 11);
  assign w271[18] = |(datain[239:236] ^ 5);
  assign w271[19] = |(datain[235:232] ^ 5);
  assign w271[20] = |(datain[231:228] ^ 7);
  assign w271[21] = |(datain[227:224] ^ 4);
  assign w271[22] = |(datain[223:220] ^ 3);
  assign w271[23] = |(datain[219:216] ^ 11);
  assign w271[24] = |(datain[215:212] ^ 2);
  assign w271[25] = |(datain[211:208] ^ 14);
  assign w271[26] = |(datain[207:204] ^ 8);
  assign w271[27] = |(datain[203:200] ^ 9);
  assign w271[28] = |(datain[199:196] ^ 8);
  assign w271[29] = |(datain[195:192] ^ 13);
  assign w271[30] = |(datain[191:188] ^ 0);
  assign w271[31] = |(datain[187:184] ^ 12);
  assign w271[32] = |(datain[183:180] ^ 0);
  assign w271[33] = |(datain[179:176] ^ 0);
  assign w271[34] = |(datain[175:172] ^ 2);
  assign w271[35] = |(datain[171:168] ^ 14);
  assign w271[36] = |(datain[167:164] ^ 8);
  assign w271[37] = |(datain[163:160] ^ 9);
  assign w271[38] = |(datain[159:156] ^ 9);
  assign w271[39] = |(datain[155:152] ^ 13);
  assign w271[40] = |(datain[151:148] ^ 0);
  assign w271[41] = |(datain[147:144] ^ 10);
  assign comp[271] = ~(|w271);
  wire [44-1:0] w272;
  assign w272[0] = |(datain[311:308] ^ 4);
  assign w272[1] = |(datain[307:304] ^ 11);
  assign w272[2] = |(datain[303:300] ^ 7);
  assign w272[3] = |(datain[299:296] ^ 5);
  assign w272[4] = |(datain[295:292] ^ 6);
  assign w272[5] = |(datain[291:288] ^ 1);
  assign w272[6] = |(datain[287:284] ^ 2);
  assign w272[7] = |(datain[283:280] ^ 14);
  assign w272[8] = |(datain[279:276] ^ 8);
  assign w272[9] = |(datain[275:272] ^ 12);
  assign w272[10] = |(datain[271:268] ^ 1);
  assign w272[11] = |(datain[267:264] ^ 14);
  assign w272[12] = |(datain[263:260] ^ 12);
  assign w272[13] = |(datain[259:256] ^ 5);
  assign w272[14] = |(datain[255:252] ^ 0);
  assign w272[15] = |(datain[251:248] ^ 1);
  assign w272[16] = |(datain[247:244] ^ 2);
  assign w272[17] = |(datain[243:240] ^ 14);
  assign w272[18] = |(datain[239:236] ^ 8);
  assign w272[19] = |(datain[235:232] ^ 9);
  assign w272[20] = |(datain[231:228] ^ 1);
  assign w272[21] = |(datain[227:224] ^ 6);
  assign w272[22] = |(datain[223:220] ^ 12);
  assign w272[23] = |(datain[219:216] ^ 7);
  assign w272[24] = |(datain[215:212] ^ 0);
  assign w272[25] = |(datain[211:208] ^ 1);
  assign w272[26] = |(datain[207:204] ^ 3);
  assign w272[27] = |(datain[203:200] ^ 2);
  assign w272[28] = |(datain[199:196] ^ 12);
  assign w272[29] = |(datain[195:192] ^ 0);
  assign w272[30] = |(datain[191:188] ^ 14);
  assign w272[31] = |(datain[187:184] ^ 8);
  assign w272[32] = |(datain[183:180] ^ 11);
  assign w272[33] = |(datain[179:176] ^ 9);
  assign w272[34] = |(datain[175:172] ^ 0);
  assign w272[35] = |(datain[171:168] ^ 2);
  assign w272[36] = |(datain[167:164] ^ 2);
  assign w272[37] = |(datain[163:160] ^ 14);
  assign w272[38] = |(datain[159:156] ^ 8);
  assign w272[39] = |(datain[155:152] ^ 9);
  assign w272[40] = |(datain[151:148] ^ 0);
  assign w272[41] = |(datain[147:144] ^ 14);
  assign w272[42] = |(datain[143:140] ^ 12);
  assign w272[43] = |(datain[139:136] ^ 9);
  assign comp[272] = ~(|w272);
  wire [44-1:0] w273;
  assign w273[0] = |(datain[311:308] ^ 1);
  assign w273[1] = |(datain[307:304] ^ 7);
  assign w273[2] = |(datain[303:300] ^ 4);
  assign w273[3] = |(datain[299:296] ^ 3);
  assign w273[4] = |(datain[295:292] ^ 3);
  assign w273[5] = |(datain[291:288] ^ 13);
  assign w273[6] = |(datain[287:284] ^ 4);
  assign w273[7] = |(datain[283:280] ^ 8);
  assign w273[8] = |(datain[279:276] ^ 0);
  assign w273[9] = |(datain[275:272] ^ 9);
  assign w273[10] = |(datain[271:268] ^ 7);
  assign w273[11] = |(datain[267:264] ^ 7);
  assign w273[12] = |(datain[263:260] ^ 0);
  assign w273[13] = |(datain[259:256] ^ 3);
  assign w273[14] = |(datain[255:252] ^ 14);
  assign w273[15] = |(datain[251:248] ^ 9);
  assign w273[16] = |(datain[247:244] ^ 0);
  assign w273[17] = |(datain[243:240] ^ 10);
  assign w273[18] = |(datain[239:236] ^ 15);
  assign w273[19] = |(datain[235:232] ^ 14);
  assign w273[20] = |(datain[231:228] ^ 3);
  assign w273[21] = |(datain[227:224] ^ 3);
  assign w273[22] = |(datain[223:220] ^ 13);
  assign w273[23] = |(datain[219:216] ^ 2);
  assign w273[24] = |(datain[215:212] ^ 9);
  assign w273[25] = |(datain[211:208] ^ 12);
  assign w273[26] = |(datain[207:204] ^ 1);
  assign w273[27] = |(datain[203:200] ^ 14);
  assign w273[28] = |(datain[199:196] ^ 5);
  assign w273[29] = |(datain[195:192] ^ 2);
  assign w273[30] = |(datain[191:188] ^ 8);
  assign w273[31] = |(datain[187:184] ^ 12);
  assign w273[32] = |(datain[183:180] ^ 12);
  assign w273[33] = |(datain[179:176] ^ 0);
  assign w273[34] = |(datain[175:172] ^ 8);
  assign w273[35] = |(datain[171:168] ^ 14);
  assign w273[36] = |(datain[167:164] ^ 13);
  assign w273[37] = |(datain[163:160] ^ 8);
  assign w273[38] = |(datain[159:156] ^ 3);
  assign w273[39] = |(datain[155:152] ^ 3);
  assign w273[40] = |(datain[151:148] ^ 12);
  assign w273[41] = |(datain[147:144] ^ 0);
  assign w273[42] = |(datain[143:140] ^ 12);
  assign w273[43] = |(datain[139:136] ^ 15);
  assign comp[273] = ~(|w273);
  wire [76-1:0] w274;
  assign w274[0] = |(datain[311:308] ^ 5);
  assign w274[1] = |(datain[307:304] ^ 0);
  assign w274[2] = |(datain[303:300] ^ 9);
  assign w274[3] = |(datain[299:296] ^ 13);
  assign w274[4] = |(datain[295:292] ^ 8);
  assign w274[5] = |(datain[291:288] ^ 11);
  assign w274[6] = |(datain[287:284] ^ 4);
  assign w274[7] = |(datain[283:280] ^ 13);
  assign w274[8] = |(datain[279:276] ^ 15);
  assign w274[9] = |(datain[275:272] ^ 12);
  assign w274[10] = |(datain[271:268] ^ 8);
  assign w274[11] = |(datain[267:264] ^ 11);
  assign w274[12] = |(datain[263:260] ^ 4);
  assign w274[13] = |(datain[259:256] ^ 5);
  assign w274[14] = |(datain[255:252] ^ 15);
  assign w274[15] = |(datain[251:248] ^ 14);
  assign w274[16] = |(datain[247:244] ^ 8);
  assign w274[17] = |(datain[243:240] ^ 10);
  assign w274[18] = |(datain[239:236] ^ 2);
  assign w274[19] = |(datain[235:232] ^ 5);
  assign w274[20] = |(datain[231:228] ^ 3);
  assign w274[21] = |(datain[227:224] ^ 2);
  assign w274[22] = |(datain[223:220] ^ 12);
  assign w274[23] = |(datain[219:216] ^ 4);
  assign w274[24] = |(datain[215:212] ^ 10);
  assign w274[25] = |(datain[211:208] ^ 10);
  assign w274[26] = |(datain[207:204] ^ 8);
  assign w274[27] = |(datain[203:200] ^ 10);
  assign w274[28] = |(datain[199:196] ^ 12);
  assign w274[29] = |(datain[195:192] ^ 4);
  assign w274[30] = |(datain[191:188] ^ 14);
  assign w274[31] = |(datain[187:184] ^ 2);
  assign w274[32] = |(datain[183:180] ^ 15);
  assign w274[33] = |(datain[179:176] ^ 7);
  assign w274[34] = |(datain[175:172] ^ 12);
  assign w274[35] = |(datain[171:168] ^ 3);
  assign w274[36] = |(datain[167:164] ^ 3);
  assign w274[37] = |(datain[163:160] ^ 3);
  assign w274[38] = |(datain[159:156] ^ 12);
  assign w274[39] = |(datain[155:152] ^ 0);
  assign w274[40] = |(datain[151:148] ^ 5);
  assign w274[41] = |(datain[147:144] ^ 0);
  assign w274[42] = |(datain[143:140] ^ 9);
  assign w274[43] = |(datain[139:136] ^ 13);
  assign w274[44] = |(datain[135:132] ^ 8);
  assign w274[45] = |(datain[131:128] ^ 11);
  assign w274[46] = |(datain[127:124] ^ 4);
  assign w274[47] = |(datain[123:120] ^ 13);
  assign w274[48] = |(datain[119:116] ^ 15);
  assign w274[49] = |(datain[115:112] ^ 12);
  assign w274[50] = |(datain[111:108] ^ 8);
  assign w274[51] = |(datain[107:104] ^ 11);
  assign w274[52] = |(datain[103:100] ^ 4);
  assign w274[53] = |(datain[99:96] ^ 5);
  assign w274[54] = |(datain[95:92] ^ 15);
  assign w274[55] = |(datain[91:88] ^ 14);
  assign w274[56] = |(datain[87:84] ^ 0);
  assign w274[57] = |(datain[83:80] ^ 2);
  assign w274[58] = |(datain[79:76] ^ 12);
  assign w274[59] = |(datain[75:72] ^ 4);
  assign w274[60] = |(datain[71:68] ^ 8);
  assign w274[61] = |(datain[67:64] ^ 9);
  assign w274[62] = |(datain[63:60] ^ 4);
  assign w274[63] = |(datain[59:56] ^ 5);
  assign w274[64] = |(datain[55:52] ^ 15);
  assign w274[65] = |(datain[51:48] ^ 14);
  assign w274[66] = |(datain[47:44] ^ 8);
  assign w274[67] = |(datain[43:40] ^ 10);
  assign w274[68] = |(datain[39:36] ^ 2);
  assign w274[69] = |(datain[35:32] ^ 5);
  assign w274[70] = |(datain[31:28] ^ 3);
  assign w274[71] = |(datain[27:24] ^ 2);
  assign w274[72] = |(datain[23:20] ^ 12);
  assign w274[73] = |(datain[19:16] ^ 4);
  assign w274[74] = |(datain[15:12] ^ 10);
  assign w274[75] = |(datain[11:8] ^ 10);
  assign comp[274] = ~(|w274);
  wire [44-1:0] w275;
  assign w275[0] = |(datain[311:308] ^ 11);
  assign w275[1] = |(datain[307:304] ^ 4);
  assign w275[2] = |(datain[303:300] ^ 3);
  assign w275[3] = |(datain[299:296] ^ 12);
  assign w275[4] = |(datain[295:292] ^ 3);
  assign w275[5] = |(datain[291:288] ^ 3);
  assign w275[6] = |(datain[287:284] ^ 12);
  assign w275[7] = |(datain[283:280] ^ 9);
  assign w275[8] = |(datain[279:276] ^ 11);
  assign w275[9] = |(datain[275:272] ^ 10);
  assign w275[10] = |(datain[271:268] ^ 9);
  assign w275[11] = |(datain[267:264] ^ 14);
  assign w275[12] = |(datain[263:260] ^ 0);
  assign w275[13] = |(datain[259:256] ^ 0);
  assign w275[14] = |(datain[255:252] ^ 12);
  assign w275[15] = |(datain[251:248] ^ 13);
  assign w275[16] = |(datain[247:244] ^ 2);
  assign w275[17] = |(datain[243:240] ^ 1);
  assign w275[18] = |(datain[239:236] ^ 11);
  assign w275[19] = |(datain[235:232] ^ 7);
  assign w275[20] = |(datain[231:228] ^ 4);
  assign w275[21] = |(datain[227:224] ^ 0);
  assign w275[22] = |(datain[223:220] ^ 9);
  assign w275[23] = |(datain[219:216] ^ 3);
  assign w275[24] = |(datain[215:212] ^ 11);
  assign w275[25] = |(datain[211:208] ^ 10);
  assign w275[26] = |(datain[207:204] ^ 0);
  assign w275[27] = |(datain[203:200] ^ 0);
  assign w275[28] = |(datain[199:196] ^ 0);
  assign w275[29] = |(datain[195:192] ^ 1);
  assign w275[30] = |(datain[191:188] ^ 11);
  assign w275[31] = |(datain[187:184] ^ 9);
  assign w275[32] = |(datain[183:180] ^ 9);
  assign w275[33] = |(datain[179:176] ^ 3);
  assign w275[34] = |(datain[175:172] ^ 0);
  assign w275[35] = |(datain[171:168] ^ 4);
  assign w275[36] = |(datain[167:164] ^ 12);
  assign w275[37] = |(datain[163:160] ^ 13);
  assign w275[38] = |(datain[159:156] ^ 2);
  assign w275[39] = |(datain[155:152] ^ 1);
  assign w275[40] = |(datain[151:148] ^ 12);
  assign w275[41] = |(datain[147:144] ^ 3);
  assign w275[42] = |(datain[143:140] ^ 11);
  assign w275[43] = |(datain[139:136] ^ 4);
  assign comp[275] = ~(|w275);
  wire [42-1:0] w276;
  assign w276[0] = |(datain[311:308] ^ 3);
  assign w276[1] = |(datain[307:304] ^ 12);
  assign w276[2] = |(datain[303:300] ^ 3);
  assign w276[3] = |(datain[299:296] ^ 3);
  assign w276[4] = |(datain[295:292] ^ 12);
  assign w276[5] = |(datain[291:288] ^ 9);
  assign w276[6] = |(datain[287:284] ^ 11);
  assign w276[7] = |(datain[283:280] ^ 10);
  assign w276[8] = |(datain[279:276] ^ 9);
  assign w276[9] = |(datain[275:272] ^ 14);
  assign w276[10] = |(datain[271:268] ^ 0);
  assign w276[11] = |(datain[267:264] ^ 0);
  assign w276[12] = |(datain[263:260] ^ 12);
  assign w276[13] = |(datain[259:256] ^ 13);
  assign w276[14] = |(datain[255:252] ^ 2);
  assign w276[15] = |(datain[251:248] ^ 1);
  assign w276[16] = |(datain[247:244] ^ 11);
  assign w276[17] = |(datain[243:240] ^ 7);
  assign w276[18] = |(datain[239:236] ^ 4);
  assign w276[19] = |(datain[235:232] ^ 0);
  assign w276[20] = |(datain[231:228] ^ 9);
  assign w276[21] = |(datain[227:224] ^ 3);
  assign w276[22] = |(datain[223:220] ^ 11);
  assign w276[23] = |(datain[219:216] ^ 10);
  assign w276[24] = |(datain[215:212] ^ 0);
  assign w276[25] = |(datain[211:208] ^ 0);
  assign w276[26] = |(datain[207:204] ^ 0);
  assign w276[27] = |(datain[203:200] ^ 1);
  assign w276[28] = |(datain[199:196] ^ 11);
  assign w276[29] = |(datain[195:192] ^ 9);
  assign w276[30] = |(datain[191:188] ^ 11);
  assign w276[31] = |(datain[187:184] ^ 0);
  assign w276[32] = |(datain[183:180] ^ 0);
  assign w276[33] = |(datain[179:176] ^ 4);
  assign w276[34] = |(datain[175:172] ^ 12);
  assign w276[35] = |(datain[171:168] ^ 13);
  assign w276[36] = |(datain[167:164] ^ 2);
  assign w276[37] = |(datain[163:160] ^ 1);
  assign w276[38] = |(datain[159:156] ^ 12);
  assign w276[39] = |(datain[155:152] ^ 3);
  assign w276[40] = |(datain[151:148] ^ 11);
  assign w276[41] = |(datain[147:144] ^ 4);
  assign comp[276] = ~(|w276);
  wire [44-1:0] w277;
  assign w277[0] = |(datain[311:308] ^ 11);
  assign w277[1] = |(datain[307:304] ^ 4);
  assign w277[2] = |(datain[303:300] ^ 3);
  assign w277[3] = |(datain[299:296] ^ 12);
  assign w277[4] = |(datain[295:292] ^ 3);
  assign w277[5] = |(datain[291:288] ^ 3);
  assign w277[6] = |(datain[287:284] ^ 12);
  assign w277[7] = |(datain[283:280] ^ 9);
  assign w277[8] = |(datain[279:276] ^ 11);
  assign w277[9] = |(datain[275:272] ^ 10);
  assign w277[10] = |(datain[271:268] ^ 9);
  assign w277[11] = |(datain[267:264] ^ 14);
  assign w277[12] = |(datain[263:260] ^ 0);
  assign w277[13] = |(datain[259:256] ^ 0);
  assign w277[14] = |(datain[255:252] ^ 12);
  assign w277[15] = |(datain[251:248] ^ 13);
  assign w277[16] = |(datain[247:244] ^ 2);
  assign w277[17] = |(datain[243:240] ^ 1);
  assign w277[18] = |(datain[239:236] ^ 11);
  assign w277[19] = |(datain[235:232] ^ 7);
  assign w277[20] = |(datain[231:228] ^ 4);
  assign w277[21] = |(datain[227:224] ^ 0);
  assign w277[22] = |(datain[223:220] ^ 9);
  assign w277[23] = |(datain[219:216] ^ 3);
  assign w277[24] = |(datain[215:212] ^ 11);
  assign w277[25] = |(datain[211:208] ^ 10);
  assign w277[26] = |(datain[207:204] ^ 0);
  assign w277[27] = |(datain[203:200] ^ 0);
  assign w277[28] = |(datain[199:196] ^ 0);
  assign w277[29] = |(datain[195:192] ^ 1);
  assign w277[30] = |(datain[191:188] ^ 11);
  assign w277[31] = |(datain[187:184] ^ 9);
  assign w277[32] = |(datain[183:180] ^ 11);
  assign w277[33] = |(datain[179:176] ^ 14);
  assign w277[34] = |(datain[175:172] ^ 0);
  assign w277[35] = |(datain[171:168] ^ 4);
  assign w277[36] = |(datain[167:164] ^ 12);
  assign w277[37] = |(datain[163:160] ^ 13);
  assign w277[38] = |(datain[159:156] ^ 2);
  assign w277[39] = |(datain[155:152] ^ 1);
  assign w277[40] = |(datain[151:148] ^ 12);
  assign w277[41] = |(datain[147:144] ^ 3);
  assign w277[42] = |(datain[143:140] ^ 11);
  assign w277[43] = |(datain[139:136] ^ 4);
  assign comp[277] = ~(|w277);
  wire [44-1:0] w278;
  assign w278[0] = |(datain[311:308] ^ 8);
  assign w278[1] = |(datain[307:304] ^ 14);
  assign w278[2] = |(datain[303:300] ^ 12);
  assign w278[3] = |(datain[299:296] ^ 0);
  assign w278[4] = |(datain[295:292] ^ 2);
  assign w278[5] = |(datain[291:288] ^ 6);
  assign w278[6] = |(datain[287:284] ^ 8);
  assign w278[7] = |(datain[283:280] ^ 3);
  assign w278[8] = |(datain[279:276] ^ 3);
  assign w278[9] = |(datain[275:272] ^ 14);
  assign w278[10] = |(datain[271:268] ^ 1);
  assign w278[11] = |(datain[267:264] ^ 8);
  assign w278[12] = |(datain[263:260] ^ 0);
  assign w278[13] = |(datain[259:256] ^ 2);
  assign w278[14] = |(datain[255:252] ^ 4);
  assign w278[15] = |(datain[251:248] ^ 0);
  assign w278[16] = |(datain[247:244] ^ 7);
  assign w278[17] = |(datain[243:240] ^ 4);
  assign w278[18] = |(datain[239:236] ^ 2);
  assign w278[19] = |(datain[235:232] ^ 10);
  assign w278[20] = |(datain[231:228] ^ 2);
  assign w278[21] = |(datain[227:224] ^ 6);
  assign w278[22] = |(datain[223:220] ^ 12);
  assign w278[23] = |(datain[219:216] ^ 7);
  assign w278[24] = |(datain[215:212] ^ 0);
  assign w278[25] = |(datain[211:208] ^ 6);
  assign w278[26] = |(datain[207:204] ^ 1);
  assign w278[27] = |(datain[203:200] ^ 8);
  assign w278[28] = |(datain[199:196] ^ 0);
  assign w278[29] = |(datain[195:192] ^ 2);
  assign w278[30] = |(datain[191:188] ^ 4);
  assign w278[31] = |(datain[187:184] ^ 0);
  assign w278[32] = |(datain[183:180] ^ 0);
  assign w278[33] = |(datain[179:176] ^ 0);
  assign w278[34] = |(datain[175:172] ^ 2);
  assign w278[35] = |(datain[171:168] ^ 6);
  assign w278[36] = |(datain[167:164] ^ 10);
  assign w278[37] = |(datain[163:160] ^ 1);
  assign w278[38] = |(datain[159:156] ^ 2);
  assign w278[39] = |(datain[155:152] ^ 0);
  assign w278[40] = |(datain[151:148] ^ 0);
  assign w278[41] = |(datain[147:144] ^ 0);
  assign w278[42] = |(datain[143:140] ^ 2);
  assign w278[43] = |(datain[139:136] ^ 6);
  assign comp[278] = ~(|w278);
  wire [46-1:0] w279;
  assign w279[0] = |(datain[311:308] ^ 0);
  assign w279[1] = |(datain[307:304] ^ 2);
  assign w279[2] = |(datain[303:300] ^ 0);
  assign w279[3] = |(datain[299:296] ^ 0);
  assign w279[4] = |(datain[295:292] ^ 11);
  assign w279[5] = |(datain[291:288] ^ 4);
  assign w279[6] = |(datain[287:284] ^ 4);
  assign w279[7] = |(datain[283:280] ^ 14);
  assign w279[8] = |(datain[279:276] ^ 11);
  assign w279[9] = |(datain[275:272] ^ 10);
  assign w279[10] = |(datain[271:268] ^ 10);
  assign w279[11] = |(datain[267:264] ^ 8);
  assign w279[12] = |(datain[263:260] ^ 0);
  assign w279[13] = |(datain[259:256] ^ 1);
  assign w279[14] = |(datain[255:252] ^ 9);
  assign w279[15] = |(datain[251:248] ^ 0);
  assign w279[16] = |(datain[247:244] ^ 12);
  assign w279[17] = |(datain[243:240] ^ 13);
  assign w279[18] = |(datain[239:236] ^ 2);
  assign w279[19] = |(datain[235:232] ^ 1);
  assign w279[20] = |(datain[231:228] ^ 11);
  assign w279[21] = |(datain[227:224] ^ 8);
  assign w279[22] = |(datain[223:220] ^ 0);
  assign w279[23] = |(datain[219:216] ^ 2);
  assign w279[24] = |(datain[215:212] ^ 3);
  assign w279[25] = |(datain[211:208] ^ 12);
  assign w279[26] = |(datain[207:204] ^ 3);
  assign w279[27] = |(datain[203:200] ^ 3);
  assign w279[28] = |(datain[199:196] ^ 12);
  assign w279[29] = |(datain[195:192] ^ 9);
  assign w279[30] = |(datain[191:188] ^ 11);
  assign w279[31] = |(datain[187:184] ^ 10);
  assign w279[32] = |(datain[183:180] ^ 9);
  assign w279[33] = |(datain[179:176] ^ 14);
  assign w279[34] = |(datain[175:172] ^ 0);
  assign w279[35] = |(datain[171:168] ^ 0);
  assign w279[36] = |(datain[167:164] ^ 12);
  assign w279[37] = |(datain[163:160] ^ 13);
  assign w279[38] = |(datain[159:156] ^ 2);
  assign w279[39] = |(datain[155:152] ^ 1);
  assign w279[40] = |(datain[151:148] ^ 11);
  assign w279[41] = |(datain[147:144] ^ 7);
  assign w279[42] = |(datain[143:140] ^ 4);
  assign w279[43] = |(datain[139:136] ^ 0);
  assign w279[44] = |(datain[135:132] ^ 9);
  assign w279[45] = |(datain[131:128] ^ 3);
  assign comp[279] = ~(|w279);
  wire [44-1:0] w280;
  assign w280[0] = |(datain[311:308] ^ 11);
  assign w280[1] = |(datain[307:304] ^ 4);
  assign w280[2] = |(datain[303:300] ^ 3);
  assign w280[3] = |(datain[299:296] ^ 12);
  assign w280[4] = |(datain[295:292] ^ 3);
  assign w280[5] = |(datain[291:288] ^ 3);
  assign w280[6] = |(datain[287:284] ^ 12);
  assign w280[7] = |(datain[283:280] ^ 9);
  assign w280[8] = |(datain[279:276] ^ 11);
  assign w280[9] = |(datain[275:272] ^ 10);
  assign w280[10] = |(datain[271:268] ^ 9);
  assign w280[11] = |(datain[267:264] ^ 14);
  assign w280[12] = |(datain[263:260] ^ 0);
  assign w280[13] = |(datain[259:256] ^ 0);
  assign w280[14] = |(datain[255:252] ^ 12);
  assign w280[15] = |(datain[251:248] ^ 13);
  assign w280[16] = |(datain[247:244] ^ 2);
  assign w280[17] = |(datain[243:240] ^ 1);
  assign w280[18] = |(datain[239:236] ^ 11);
  assign w280[19] = |(datain[235:232] ^ 7);
  assign w280[20] = |(datain[231:228] ^ 4);
  assign w280[21] = |(datain[227:224] ^ 0);
  assign w280[22] = |(datain[223:220] ^ 9);
  assign w280[23] = |(datain[219:216] ^ 3);
  assign w280[24] = |(datain[215:212] ^ 11);
  assign w280[25] = |(datain[211:208] ^ 10);
  assign w280[26] = |(datain[207:204] ^ 0);
  assign w280[27] = |(datain[203:200] ^ 0);
  assign w280[28] = |(datain[199:196] ^ 0);
  assign w280[29] = |(datain[195:192] ^ 1);
  assign w280[30] = |(datain[191:188] ^ 11);
  assign w280[31] = |(datain[187:184] ^ 9);
  assign w280[32] = |(datain[183:180] ^ 9);
  assign w280[33] = |(datain[179:176] ^ 2);
  assign w280[34] = |(datain[175:172] ^ 0);
  assign w280[35] = |(datain[171:168] ^ 4);
  assign w280[36] = |(datain[167:164] ^ 12);
  assign w280[37] = |(datain[163:160] ^ 13);
  assign w280[38] = |(datain[159:156] ^ 2);
  assign w280[39] = |(datain[155:152] ^ 1);
  assign w280[40] = |(datain[151:148] ^ 12);
  assign w280[41] = |(datain[147:144] ^ 3);
  assign w280[42] = |(datain[143:140] ^ 11);
  assign w280[43] = |(datain[139:136] ^ 4);
  assign comp[280] = ~(|w280);
  wire [56-1:0] w281;
  assign w281[0] = |(datain[311:308] ^ 3);
  assign w281[1] = |(datain[307:304] ^ 12);
  assign w281[2] = |(datain[303:300] ^ 3);
  assign w281[3] = |(datain[299:296] ^ 3);
  assign w281[4] = |(datain[295:292] ^ 12);
  assign w281[5] = |(datain[291:288] ^ 9);
  assign w281[6] = |(datain[287:284] ^ 11);
  assign w281[7] = |(datain[283:280] ^ 10);
  assign w281[8] = |(datain[279:276] ^ 9);
  assign w281[9] = |(datain[275:272] ^ 14);
  assign w281[10] = |(datain[271:268] ^ 0);
  assign w281[11] = |(datain[267:264] ^ 0);
  assign w281[12] = |(datain[263:260] ^ 12);
  assign w281[13] = |(datain[259:256] ^ 13);
  assign w281[14] = |(datain[255:252] ^ 2);
  assign w281[15] = |(datain[251:248] ^ 1);
  assign w281[16] = |(datain[247:244] ^ 11);
  assign w281[17] = |(datain[243:240] ^ 7);
  assign w281[18] = |(datain[239:236] ^ 4);
  assign w281[19] = |(datain[235:232] ^ 0);
  assign w281[20] = |(datain[231:228] ^ 9);
  assign w281[21] = |(datain[227:224] ^ 3);
  assign w281[22] = |(datain[223:220] ^ 11);
  assign w281[23] = |(datain[219:216] ^ 10);
  assign w281[24] = |(datain[215:212] ^ 0);
  assign w281[25] = |(datain[211:208] ^ 0);
  assign w281[26] = |(datain[207:204] ^ 0);
  assign w281[27] = |(datain[203:200] ^ 1);
  assign w281[28] = |(datain[199:196] ^ 11);
  assign w281[29] = |(datain[195:192] ^ 9);
  assign w281[30] = |(datain[191:188] ^ 12);
  assign w281[31] = |(datain[187:184] ^ 3);
  assign w281[32] = |(datain[183:180] ^ 0);
  assign w281[33] = |(datain[179:176] ^ 4);
  assign w281[34] = |(datain[175:172] ^ 12);
  assign w281[35] = |(datain[171:168] ^ 13);
  assign w281[36] = |(datain[167:164] ^ 2);
  assign w281[37] = |(datain[163:160] ^ 1);
  assign w281[38] = |(datain[159:156] ^ 12);
  assign w281[39] = |(datain[155:152] ^ 3);
  assign w281[40] = |(datain[151:148] ^ 11);
  assign w281[41] = |(datain[147:144] ^ 4);
  assign w281[42] = |(datain[143:140] ^ 3);
  assign w281[43] = |(datain[139:136] ^ 11);
  assign w281[44] = |(datain[135:132] ^ 11);
  assign w281[45] = |(datain[131:128] ^ 10);
  assign w281[46] = |(datain[127:124] ^ 11);
  assign w281[47] = |(datain[123:120] ^ 14);
  assign w281[48] = |(datain[119:116] ^ 0);
  assign w281[49] = |(datain[115:112] ^ 1);
  assign w281[50] = |(datain[111:108] ^ 12);
  assign w281[51] = |(datain[107:104] ^ 13);
  assign w281[52] = |(datain[103:100] ^ 2);
  assign w281[53] = |(datain[99:96] ^ 1);
  assign w281[54] = |(datain[95:92] ^ 12);
  assign w281[55] = |(datain[91:88] ^ 3);
  assign comp[281] = ~(|w281);
  wire [76-1:0] w282;
  assign w282[0] = |(datain[311:308] ^ 4);
  assign w282[1] = |(datain[307:304] ^ 4);
  assign w282[2] = |(datain[303:300] ^ 15);
  assign w282[3] = |(datain[299:296] ^ 13);
  assign w282[4] = |(datain[295:292] ^ 14);
  assign w282[5] = |(datain[291:288] ^ 9);
  assign w282[6] = |(datain[287:284] ^ 8);
  assign w282[7] = |(datain[283:280] ^ 9);
  assign w282[8] = |(datain[279:276] ^ 4);
  assign w282[9] = |(datain[275:272] ^ 4);
  assign w282[10] = |(datain[271:268] ^ 15);
  assign w282[11] = |(datain[267:264] ^ 14);
  assign w282[12] = |(datain[263:260] ^ 11);
  assign w282[13] = |(datain[259:256] ^ 4);
  assign w282[14] = |(datain[255:252] ^ 4);
  assign w282[15] = |(datain[251:248] ^ 0);
  assign w282[16] = |(datain[247:244] ^ 8);
  assign w282[17] = |(datain[243:240] ^ 13);
  assign w282[18] = |(datain[239:236] ^ 9);
  assign w282[19] = |(datain[235:232] ^ 6);
  assign w282[20] = |(datain[231:228] ^ 0);
  assign w282[21] = |(datain[227:224] ^ 3);
  assign w282[22] = |(datain[223:220] ^ 0);
  assign w282[23] = |(datain[219:216] ^ 1);
  assign w282[24] = |(datain[215:212] ^ 11);
  assign w282[25] = |(datain[211:208] ^ 9);
  assign w282[26] = |(datain[207:204] ^ 13);
  assign w282[27] = |(datain[203:200] ^ 11);
  assign w282[28] = |(datain[199:196] ^ 0);
  assign w282[29] = |(datain[195:192] ^ 7);
  assign w282[30] = |(datain[191:188] ^ 12);
  assign w282[31] = |(datain[187:184] ^ 13);
  assign w282[32] = |(datain[183:180] ^ 2);
  assign w282[33] = |(datain[179:176] ^ 1);
  assign w282[34] = |(datain[175:172] ^ 11);
  assign w282[35] = |(datain[171:168] ^ 8);
  assign w282[36] = |(datain[167:164] ^ 0);
  assign w282[37] = |(datain[163:160] ^ 0);
  assign w282[38] = |(datain[159:156] ^ 4);
  assign w282[39] = |(datain[155:152] ^ 2);
  assign w282[40] = |(datain[151:148] ^ 3);
  assign w282[41] = |(datain[147:144] ^ 3);
  assign w282[42] = |(datain[143:140] ^ 12);
  assign w282[43] = |(datain[139:136] ^ 9);
  assign w282[44] = |(datain[135:132] ^ 9);
  assign w282[45] = |(datain[131:128] ^ 9);
  assign w282[46] = |(datain[127:124] ^ 12);
  assign w282[47] = |(datain[123:120] ^ 13);
  assign w282[48] = |(datain[119:116] ^ 2);
  assign w282[49] = |(datain[115:112] ^ 1);
  assign w282[50] = |(datain[111:108] ^ 11);
  assign w282[51] = |(datain[107:104] ^ 4);
  assign w282[52] = |(datain[103:100] ^ 4);
  assign w282[53] = |(datain[99:96] ^ 0);
  assign w282[54] = |(datain[95:92] ^ 8);
  assign w282[55] = |(datain[91:88] ^ 13);
  assign w282[56] = |(datain[87:84] ^ 9);
  assign w282[57] = |(datain[83:80] ^ 6);
  assign w282[58] = |(datain[79:76] ^ 4);
  assign w282[59] = |(datain[75:72] ^ 11);
  assign w282[60] = |(datain[71:68] ^ 0);
  assign w282[61] = |(datain[67:64] ^ 9);
  assign w282[62] = |(datain[63:60] ^ 5);
  assign w282[63] = |(datain[59:56] ^ 9);
  assign w282[64] = |(datain[55:52] ^ 12);
  assign w282[65] = |(datain[51:48] ^ 13);
  assign w282[66] = |(datain[47:44] ^ 2);
  assign w282[67] = |(datain[43:40] ^ 1);
  assign w282[68] = |(datain[39:36] ^ 15);
  assign w282[69] = |(datain[35:32] ^ 14);
  assign w282[70] = |(datain[31:28] ^ 8);
  assign w282[71] = |(datain[27:24] ^ 14);
  assign w282[72] = |(datain[23:20] ^ 4);
  assign w282[73] = |(datain[19:16] ^ 10);
  assign w282[74] = |(datain[15:12] ^ 0);
  assign w282[75] = |(datain[11:8] ^ 9);
  assign comp[282] = ~(|w282);
  wire [74-1:0] w283;
  assign w283[0] = |(datain[311:308] ^ 11);
  assign w283[1] = |(datain[307:304] ^ 4);
  assign w283[2] = |(datain[303:300] ^ 3);
  assign w283[3] = |(datain[299:296] ^ 13);
  assign w283[4] = |(datain[295:292] ^ 8);
  assign w283[5] = |(datain[291:288] ^ 13);
  assign w283[6] = |(datain[287:284] ^ 9);
  assign w283[7] = |(datain[283:280] ^ 6);
  assign w283[8] = |(datain[279:276] ^ 8);
  assign w283[9] = |(datain[275:272] ^ 4);
  assign w283[10] = |(datain[271:268] ^ 0);
  assign w283[11] = |(datain[267:264] ^ 3);
  assign w283[12] = |(datain[263:260] ^ 12);
  assign w283[13] = |(datain[259:256] ^ 13);
  assign w283[14] = |(datain[255:252] ^ 2);
  assign w283[15] = |(datain[251:248] ^ 1);
  assign w283[16] = |(datain[247:244] ^ 9);
  assign w283[17] = |(datain[243:240] ^ 3);
  assign w283[18] = |(datain[239:236] ^ 12);
  assign w283[19] = |(datain[235:232] ^ 3);
  assign w283[20] = |(datain[231:228] ^ 11);
  assign w283[21] = |(datain[227:224] ^ 8);
  assign w283[22] = |(datain[223:220] ^ 0);
  assign w283[23] = |(datain[219:216] ^ 1);
  assign w283[24] = |(datain[215:212] ^ 4);
  assign w283[25] = |(datain[211:208] ^ 3);
  assign w283[26] = |(datain[207:204] ^ 8);
  assign w283[27] = |(datain[203:200] ^ 13);
  assign w283[28] = |(datain[199:196] ^ 9);
  assign w283[29] = |(datain[195:192] ^ 6);
  assign w283[30] = |(datain[191:188] ^ 8);
  assign w283[31] = |(datain[187:184] ^ 4);
  assign w283[32] = |(datain[183:180] ^ 0);
  assign w283[33] = |(datain[179:176] ^ 3);
  assign w283[34] = |(datain[175:172] ^ 12);
  assign w283[35] = |(datain[171:168] ^ 13);
  assign w283[36] = |(datain[167:164] ^ 2);
  assign w283[37] = |(datain[163:160] ^ 1);
  assign w283[38] = |(datain[159:156] ^ 12);
  assign w283[39] = |(datain[155:152] ^ 3);
  assign w283[40] = |(datain[151:148] ^ 5);
  assign w283[41] = |(datain[147:144] ^ 11);
  assign w283[42] = |(datain[143:140] ^ 5);
  assign w283[43] = |(datain[139:136] ^ 13);
  assign w283[44] = |(datain[135:132] ^ 11);
  assign w283[45] = |(datain[131:128] ^ 4);
  assign w283[46] = |(datain[127:124] ^ 4);
  assign w283[47] = |(datain[123:120] ^ 0);
  assign w283[48] = |(datain[119:116] ^ 8);
  assign w283[49] = |(datain[115:112] ^ 13);
  assign w283[50] = |(datain[111:108] ^ 9);
  assign w283[51] = |(datain[107:104] ^ 6);
  assign w283[52] = |(datain[103:100] ^ 0);
  assign w283[53] = |(datain[99:96] ^ 3);
  assign w283[54] = |(datain[95:92] ^ 0);
  assign w283[55] = |(datain[91:88] ^ 1);
  assign w283[56] = |(datain[87:84] ^ 11);
  assign w283[57] = |(datain[83:80] ^ 9);
  assign w283[58] = |(datain[79:76] ^ 12);
  assign w283[59] = |(datain[75:72] ^ 10);
  assign w283[60] = |(datain[71:68] ^ 0);
  assign w283[61] = |(datain[67:64] ^ 1);
  assign w283[62] = |(datain[63:60] ^ 12);
  assign w283[63] = |(datain[59:56] ^ 13);
  assign w283[64] = |(datain[55:52] ^ 2);
  assign w283[65] = |(datain[51:48] ^ 1);
  assign w283[66] = |(datain[47:44] ^ 5);
  assign w283[67] = |(datain[43:40] ^ 3);
  assign w283[68] = |(datain[39:36] ^ 5);
  assign w283[69] = |(datain[35:32] ^ 5);
  assign w283[70] = |(datain[31:28] ^ 11);
  assign w283[71] = |(datain[27:24] ^ 0);
  assign w283[72] = |(datain[23:20] ^ 0);
  assign w283[73] = |(datain[19:16] ^ 3);
  assign comp[283] = ~(|w283);
  wire [76-1:0] w284;
  assign w284[0] = |(datain[311:308] ^ 0);
  assign w284[1] = |(datain[307:304] ^ 7);
  assign w284[2] = |(datain[303:300] ^ 8);
  assign w284[3] = |(datain[299:296] ^ 14);
  assign w284[4] = |(datain[295:292] ^ 13);
  assign w284[5] = |(datain[291:288] ^ 0);
  assign w284[6] = |(datain[287:284] ^ 3);
  assign w284[7] = |(datain[283:280] ^ 3);
  assign w284[8] = |(datain[279:276] ^ 14);
  assign w284[9] = |(datain[275:272] ^ 4);
  assign w284[10] = |(datain[271:268] ^ 8);
  assign w284[11] = |(datain[267:264] ^ 14);
  assign w284[12] = |(datain[263:260] ^ 13);
  assign w284[13] = |(datain[259:256] ^ 8);
  assign w284[14] = |(datain[255:252] ^ 8);
  assign w284[15] = |(datain[251:248] ^ 14);
  assign w284[16] = |(datain[247:244] ^ 12);
  assign w284[17] = |(datain[243:240] ^ 0);
  assign w284[18] = |(datain[239:236] ^ 1);
  assign w284[19] = |(datain[235:232] ^ 14);
  assign w284[20] = |(datain[231:228] ^ 3);
  assign w284[21] = |(datain[227:224] ^ 3);
  assign w284[22] = |(datain[223:220] ^ 12);
  assign w284[23] = |(datain[219:216] ^ 0);
  assign w284[24] = |(datain[215:212] ^ 10);
  assign w284[25] = |(datain[211:208] ^ 3);
  assign w284[26] = |(datain[207:204] ^ 8);
  assign w284[27] = |(datain[203:200] ^ 1);
  assign w284[28] = |(datain[199:196] ^ 0);
  assign w284[29] = |(datain[195:192] ^ 0);
  assign w284[30] = |(datain[191:188] ^ 8);
  assign w284[31] = |(datain[187:184] ^ 14);
  assign w284[32] = |(datain[183:180] ^ 13);
  assign w284[33] = |(datain[179:176] ^ 8);
  assign w284[34] = |(datain[175:172] ^ 1);
  assign w284[35] = |(datain[171:168] ^ 14);
  assign w284[36] = |(datain[167:164] ^ 8);
  assign w284[37] = |(datain[163:160] ^ 11);
  assign w284[38] = |(datain[159:156] ^ 15);
  assign w284[39] = |(datain[155:152] ^ 0);
  assign w284[40] = |(datain[151:148] ^ 8);
  assign w284[41] = |(datain[147:144] ^ 11);
  assign w284[42] = |(datain[143:140] ^ 15);
  assign w284[43] = |(datain[139:136] ^ 8);
  assign w284[44] = |(datain[135:132] ^ 15);
  assign w284[45] = |(datain[131:128] ^ 15);
  assign w284[46] = |(datain[127:124] ^ 0);
  assign w284[47] = |(datain[123:120] ^ 14);
  assign w284[48] = |(datain[119:116] ^ 1);
  assign w284[49] = |(datain[115:112] ^ 3);
  assign w284[50] = |(datain[111:108] ^ 0);
  assign w284[51] = |(datain[107:104] ^ 4);
  assign w284[52] = |(datain[103:100] ^ 10);
  assign w284[53] = |(datain[99:96] ^ 1);
  assign w284[54] = |(datain[95:92] ^ 1);
  assign w284[55] = |(datain[91:88] ^ 3);
  assign w284[56] = |(datain[87:84] ^ 0);
  assign w284[57] = |(datain[83:80] ^ 4);
  assign w284[58] = |(datain[79:76] ^ 11);
  assign w284[59] = |(datain[75:72] ^ 1);
  assign w284[60] = |(datain[71:68] ^ 0);
  assign w284[61] = |(datain[67:64] ^ 6);
  assign w284[62] = |(datain[63:60] ^ 13);
  assign w284[63] = |(datain[59:56] ^ 3);
  assign w284[64] = |(datain[55:52] ^ 14);
  assign w284[65] = |(datain[51:48] ^ 0);
  assign w284[66] = |(datain[47:44] ^ 5);
  assign w284[67] = |(datain[43:40] ^ 0);
  assign w284[68] = |(datain[39:36] ^ 5);
  assign w284[69] = |(datain[35:32] ^ 0);
  assign w284[70] = |(datain[31:28] ^ 8);
  assign w284[71] = |(datain[27:24] ^ 11);
  assign w284[72] = |(datain[23:20] ^ 1);
  assign w284[73] = |(datain[19:16] ^ 14);
  assign w284[74] = |(datain[15:12] ^ 4);
  assign w284[75] = |(datain[11:8] ^ 14);
  assign comp[284] = ~(|w284);
  wire [76-1:0] w285;
  assign w285[0] = |(datain[311:308] ^ 4);
  assign w285[1] = |(datain[307:304] ^ 1);
  assign w285[2] = |(datain[303:300] ^ 7);
  assign w285[3] = |(datain[299:296] ^ 5);
  assign w285[4] = |(datain[295:292] ^ 2);
  assign w285[5] = |(datain[291:288] ^ 3);
  assign w285[6] = |(datain[287:284] ^ 10);
  assign w285[7] = |(datain[283:280] ^ 13);
  assign w285[8] = |(datain[279:276] ^ 3);
  assign w285[9] = |(datain[275:272] ^ 13);
  assign w285[10] = |(datain[271:268] ^ 2);
  assign w285[11] = |(datain[267:264] ^ 14);
  assign w285[12] = |(datain[263:260] ^ 4);
  assign w285[13] = |(datain[259:256] ^ 4);
  assign w285[14] = |(datain[255:252] ^ 7);
  assign w285[15] = |(datain[251:248] ^ 5);
  assign w285[16] = |(datain[247:244] ^ 1);
  assign w285[17] = |(datain[243:240] ^ 13);
  assign w285[18] = |(datain[239:236] ^ 10);
  assign w285[19] = |(datain[235:232] ^ 13);
  assign w285[20] = |(datain[231:228] ^ 3);
  assign w285[21] = |(datain[227:224] ^ 13);
  assign w285[22] = |(datain[223:220] ^ 4);
  assign w285[23] = |(datain[219:216] ^ 2);
  assign w285[24] = |(datain[215:212] ^ 4);
  assign w285[25] = |(datain[211:208] ^ 6);
  assign w285[26] = |(datain[207:204] ^ 7);
  assign w285[27] = |(datain[203:200] ^ 5);
  assign w285[28] = |(datain[199:196] ^ 1);
  assign w285[29] = |(datain[195:192] ^ 7);
  assign w285[30] = |(datain[191:188] ^ 11);
  assign w285[31] = |(datain[187:184] ^ 8);
  assign w285[32] = |(datain[183:180] ^ 0);
  assign w285[33] = |(datain[179:176] ^ 2);
  assign w285[34] = |(datain[175:172] ^ 3);
  assign w285[35] = |(datain[171:168] ^ 13);
  assign w285[36] = |(datain[167:164] ^ 14);
  assign w285[37] = |(datain[163:160] ^ 8);
  assign w285[38] = |(datain[159:156] ^ 1);
  assign w285[39] = |(datain[155:152] ^ 7);
  assign w285[40] = |(datain[151:148] ^ 0);
  assign w285[41] = |(datain[147:144] ^ 0);
  assign w285[42] = |(datain[143:140] ^ 8);
  assign w285[43] = |(datain[139:136] ^ 11);
  assign w285[44] = |(datain[135:132] ^ 13);
  assign w285[45] = |(datain[131:128] ^ 8);
  assign w285[46] = |(datain[127:124] ^ 11);
  assign w285[47] = |(datain[123:120] ^ 4);
  assign w285[48] = |(datain[119:116] ^ 4);
  assign w285[49] = |(datain[115:112] ^ 0);
  assign w285[50] = |(datain[111:108] ^ 11);
  assign w285[51] = |(datain[107:104] ^ 9);
  assign w285[52] = |(datain[103:100] ^ 0);
  assign w285[53] = |(datain[99:96] ^ 0);
  assign w285[54] = |(datain[95:92] ^ 0);
  assign w285[55] = |(datain[91:88] ^ 2);
  assign w285[56] = |(datain[87:84] ^ 3);
  assign w285[57] = |(datain[83:80] ^ 3);
  assign w285[58] = |(datain[79:76] ^ 13);
  assign w285[59] = |(datain[75:72] ^ 2);
  assign w285[60] = |(datain[71:68] ^ 14);
  assign w285[61] = |(datain[67:64] ^ 8);
  assign w285[62] = |(datain[63:60] ^ 0);
  assign w285[63] = |(datain[59:56] ^ 11);
  assign w285[64] = |(datain[55:52] ^ 0);
  assign w285[65] = |(datain[51:48] ^ 0);
  assign w285[66] = |(datain[47:44] ^ 11);
  assign w285[67] = |(datain[43:40] ^ 4);
  assign w285[68] = |(datain[39:36] ^ 3);
  assign w285[69] = |(datain[35:32] ^ 14);
  assign w285[70] = |(datain[31:28] ^ 14);
  assign w285[71] = |(datain[27:24] ^ 8);
  assign w285[72] = |(datain[23:20] ^ 0);
  assign w285[73] = |(datain[19:16] ^ 6);
  assign w285[74] = |(datain[15:12] ^ 0);
  assign w285[75] = |(datain[11:8] ^ 0);
  assign comp[285] = ~(|w285);
  wire [70-1:0] w286;
  assign w286[0] = |(datain[311:308] ^ 14);
  assign w286[1] = |(datain[307:304] ^ 8);
  assign w286[2] = |(datain[303:300] ^ 0);
  assign w286[3] = |(datain[299:296] ^ 0);
  assign w286[4] = |(datain[295:292] ^ 0);
  assign w286[5] = |(datain[291:288] ^ 0);
  assign w286[6] = |(datain[287:284] ^ 8);
  assign w286[7] = |(datain[283:280] ^ 7);
  assign w286[8] = |(datain[279:276] ^ 13);
  assign w286[9] = |(datain[275:272] ^ 11);
  assign w286[10] = |(datain[271:268] ^ 5);
  assign w286[11] = |(datain[267:264] ^ 11);
  assign w286[12] = |(datain[263:260] ^ 8);
  assign w286[13] = |(datain[259:256] ^ 1);
  assign w286[14] = |(datain[255:252] ^ 14);
  assign w286[15] = |(datain[251:248] ^ 11);
  assign w286[16] = |(datain[247:244] ^ 0);
  assign w286[17] = |(datain[243:240] ^ 3);
  assign w286[18] = |(datain[239:236] ^ 0);
  assign w286[19] = |(datain[235:232] ^ 1);
  assign w286[20] = |(datain[231:228] ^ 0);
  assign w286[21] = |(datain[227:224] ^ 14);
  assign w286[22] = |(datain[223:220] ^ 1);
  assign w286[23] = |(datain[219:216] ^ 15);
  assign w286[24] = |(datain[215:212] ^ 8);
  assign w286[25] = |(datain[211:208] ^ 10);
  assign w286[26] = |(datain[207:204] ^ 8);
  assign w286[27] = |(datain[203:200] ^ 7);
  assign w286[28] = |(datain[199:196] ^ 2);
  assign w286[29] = |(datain[195:192] ^ 3);
  assign w286[30] = |(datain[191:188] ^ 0);
  assign w286[31] = |(datain[187:184] ^ 1);
  assign w286[32] = |(datain[183:180] ^ 3);
  assign w286[33] = |(datain[179:176] ^ 3);
  assign w286[34] = |(datain[175:172] ^ 15);
  assign w286[35] = |(datain[171:168] ^ 15);
  assign w286[36] = |(datain[167:164] ^ 8);
  assign w286[37] = |(datain[163:160] ^ 7);
  assign w286[38] = |(datain[159:156] ^ 12);
  assign w286[39] = |(datain[155:152] ^ 9);
  assign w286[40] = |(datain[151:148] ^ 11);
  assign w286[41] = |(datain[147:144] ^ 9);
  assign w286[42] = |(datain[143:140] ^ 15);
  assign w286[43] = |(datain[139:136] ^ 12);
  assign w286[44] = |(datain[135:132] ^ 0);
  assign w286[45] = |(datain[131:128] ^ 13);
  assign w286[46] = |(datain[127:124] ^ 9);
  assign w286[47] = |(datain[123:120] ^ 0);
  assign w286[48] = |(datain[119:116] ^ 3);
  assign w286[49] = |(datain[115:112] ^ 0);
  assign w286[50] = |(datain[111:108] ^ 8);
  assign w286[51] = |(datain[107:104] ^ 1);
  assign w286[52] = |(datain[103:100] ^ 2);
  assign w286[53] = |(datain[99:96] ^ 7);
  assign w286[54] = |(datain[95:92] ^ 0);
  assign w286[55] = |(datain[91:88] ^ 1);
  assign w286[56] = |(datain[87:84] ^ 8);
  assign w286[57] = |(datain[83:80] ^ 7);
  assign w286[58] = |(datain[79:76] ^ 13);
  assign w286[59] = |(datain[75:72] ^ 2);
  assign w286[60] = |(datain[71:68] ^ 4);
  assign w286[61] = |(datain[67:64] ^ 7);
  assign w286[62] = |(datain[63:60] ^ 14);
  assign w286[63] = |(datain[59:56] ^ 2);
  assign w286[64] = |(datain[55:52] ^ 15);
  assign w286[65] = |(datain[51:48] ^ 7);
  assign w286[66] = |(datain[47:44] ^ 14);
  assign w286[67] = |(datain[43:40] ^ 11);
  assign w286[68] = |(datain[39:36] ^ 0);
  assign w286[69] = |(datain[35:32] ^ 4);
  assign comp[286] = ~(|w286);
  wire [64-1:0] w287;
  assign w287[0] = |(datain[311:308] ^ 8);
  assign w287[1] = |(datain[307:304] ^ 7);
  assign w287[2] = |(datain[303:300] ^ 13);
  assign w287[3] = |(datain[299:296] ^ 11);
  assign w287[4] = |(datain[295:292] ^ 5);
  assign w287[5] = |(datain[291:288] ^ 11);
  assign w287[6] = |(datain[287:284] ^ 8);
  assign w287[7] = |(datain[283:280] ^ 1);
  assign w287[8] = |(datain[279:276] ^ 14);
  assign w287[9] = |(datain[275:272] ^ 11);
  assign w287[10] = |(datain[271:268] ^ 0);
  assign w287[11] = |(datain[267:264] ^ 3);
  assign w287[12] = |(datain[263:260] ^ 0);
  assign w287[13] = |(datain[259:256] ^ 1);
  assign w287[14] = |(datain[255:252] ^ 0);
  assign w287[15] = |(datain[251:248] ^ 14);
  assign w287[16] = |(datain[247:244] ^ 1);
  assign w287[17] = |(datain[243:240] ^ 15);
  assign w287[18] = |(datain[239:236] ^ 8);
  assign w287[19] = |(datain[235:232] ^ 10);
  assign w287[20] = |(datain[231:228] ^ 8);
  assign w287[21] = |(datain[227:224] ^ 7);
  assign w287[22] = |(datain[223:220] ^ 2);
  assign w287[23] = |(datain[219:216] ^ 3);
  assign w287[24] = |(datain[215:212] ^ 0);
  assign w287[25] = |(datain[211:208] ^ 1);
  assign w287[26] = |(datain[207:204] ^ 3);
  assign w287[27] = |(datain[203:200] ^ 3);
  assign w287[28] = |(datain[199:196] ^ 15);
  assign w287[29] = |(datain[195:192] ^ 15);
  assign w287[30] = |(datain[191:188] ^ 8);
  assign w287[31] = |(datain[187:184] ^ 7);
  assign w287[32] = |(datain[183:180] ^ 12);
  assign w287[33] = |(datain[179:176] ^ 9);
  assign w287[34] = |(datain[175:172] ^ 11);
  assign w287[35] = |(datain[171:168] ^ 9);
  assign w287[36] = |(datain[167:164] ^ 9);
  assign w287[37] = |(datain[163:160] ^ 6);
  assign w287[38] = |(datain[159:156] ^ 0);
  assign w287[39] = |(datain[155:152] ^ 14);
  assign w287[40] = |(datain[151:148] ^ 9);
  assign w287[41] = |(datain[147:144] ^ 0);
  assign w287[42] = |(datain[143:140] ^ 3);
  assign w287[43] = |(datain[139:136] ^ 0);
  assign w287[44] = |(datain[135:132] ^ 8);
  assign w287[45] = |(datain[131:128] ^ 1);
  assign w287[46] = |(datain[127:124] ^ 2);
  assign w287[47] = |(datain[123:120] ^ 7);
  assign w287[48] = |(datain[119:116] ^ 0);
  assign w287[49] = |(datain[115:112] ^ 1);
  assign w287[50] = |(datain[111:108] ^ 8);
  assign w287[51] = |(datain[107:104] ^ 7);
  assign w287[52] = |(datain[103:100] ^ 13);
  assign w287[53] = |(datain[99:96] ^ 2);
  assign w287[54] = |(datain[95:92] ^ 4);
  assign w287[55] = |(datain[91:88] ^ 7);
  assign w287[56] = |(datain[87:84] ^ 14);
  assign w287[57] = |(datain[83:80] ^ 2);
  assign w287[58] = |(datain[79:76] ^ 15);
  assign w287[59] = |(datain[75:72] ^ 7);
  assign w287[60] = |(datain[71:68] ^ 14);
  assign w287[61] = |(datain[67:64] ^ 11);
  assign w287[62] = |(datain[63:60] ^ 0);
  assign w287[63] = |(datain[59:56] ^ 4);
  assign comp[287] = ~(|w287);
  wire [74-1:0] w288;
  assign w288[0] = |(datain[311:308] ^ 0);
  assign w288[1] = |(datain[307:304] ^ 3);
  assign w288[2] = |(datain[303:300] ^ 14);
  assign w288[3] = |(datain[299:296] ^ 9);
  assign w288[4] = |(datain[295:292] ^ 10);
  assign w288[5] = |(datain[291:288] ^ 1);
  assign w288[6] = |(datain[287:284] ^ 1);
  assign w288[7] = |(datain[283:280] ^ 9);
  assign w288[8] = |(datain[279:276] ^ 0);
  assign w288[9] = |(datain[275:272] ^ 3);
  assign w288[10] = |(datain[271:268] ^ 2);
  assign w288[11] = |(datain[267:264] ^ 13);
  assign w288[12] = |(datain[263:260] ^ 0);
  assign w288[13] = |(datain[259:256] ^ 3);
  assign w288[14] = |(datain[255:252] ^ 0);
  assign w288[15] = |(datain[251:248] ^ 0);
  assign w288[16] = |(datain[247:244] ^ 10);
  assign w288[17] = |(datain[243:240] ^ 3);
  assign w288[18] = |(datain[239:236] ^ 3);
  assign w288[19] = |(datain[235:232] ^ 1);
  assign w288[20] = |(datain[231:228] ^ 0);
  assign w288[21] = |(datain[227:224] ^ 3);
  assign w288[22] = |(datain[223:220] ^ 11);
  assign w288[23] = |(datain[219:216] ^ 4);
  assign w288[24] = |(datain[215:212] ^ 4);
  assign w288[25] = |(datain[211:208] ^ 0);
  assign w288[26] = |(datain[207:204] ^ 11);
  assign w288[27] = |(datain[203:200] ^ 9);
  assign w288[28] = |(datain[199:196] ^ 0);
  assign w288[29] = |(datain[195:192] ^ 3);
  assign w288[30] = |(datain[191:188] ^ 0);
  assign w288[31] = |(datain[187:184] ^ 0);
  assign w288[32] = |(datain[183:180] ^ 11);
  assign w288[33] = |(datain[179:176] ^ 10);
  assign w288[34] = |(datain[175:172] ^ 3);
  assign w288[35] = |(datain[171:168] ^ 0);
  assign w288[36] = |(datain[167:164] ^ 0);
  assign w288[37] = |(datain[163:160] ^ 3);
  assign w288[38] = |(datain[159:156] ^ 12);
  assign w288[39] = |(datain[155:152] ^ 13);
  assign w288[40] = |(datain[151:148] ^ 2);
  assign w288[41] = |(datain[147:144] ^ 1);
  assign w288[42] = |(datain[143:140] ^ 11);
  assign w288[43] = |(datain[139:136] ^ 8);
  assign w288[44] = |(datain[135:132] ^ 0);
  assign w288[45] = |(datain[131:128] ^ 1);
  assign w288[46] = |(datain[127:124] ^ 5);
  assign w288[47] = |(datain[123:120] ^ 7);
  assign w288[48] = |(datain[119:116] ^ 8);
  assign w288[49] = |(datain[115:112] ^ 11);
  assign w288[50] = |(datain[111:108] ^ 0);
  assign w288[51] = |(datain[107:104] ^ 14);
  assign w288[52] = |(datain[103:100] ^ 1);
  assign w288[53] = |(datain[99:96] ^ 5);
  assign w288[54] = |(datain[95:92] ^ 0);
  assign w288[55] = |(datain[91:88] ^ 3);
  assign w288[56] = |(datain[87:84] ^ 8);
  assign w288[57] = |(datain[83:80] ^ 0);
  assign w288[58] = |(datain[79:76] ^ 12);
  assign w288[59] = |(datain[75:72] ^ 9);
  assign w288[60] = |(datain[71:68] ^ 1);
  assign w288[61] = |(datain[67:64] ^ 15);
  assign w288[62] = |(datain[63:60] ^ 8);
  assign w288[63] = |(datain[59:56] ^ 11);
  assign w288[64] = |(datain[55:52] ^ 1);
  assign w288[65] = |(datain[51:48] ^ 6);
  assign w288[66] = |(datain[47:44] ^ 1);
  assign w288[67] = |(datain[43:40] ^ 7);
  assign w288[68] = |(datain[39:36] ^ 0);
  assign w288[69] = |(datain[35:32] ^ 3);
  assign w288[70] = |(datain[31:28] ^ 12);
  assign w288[71] = |(datain[27:24] ^ 13);
  assign w288[72] = |(datain[23:20] ^ 2);
  assign w288[73] = |(datain[19:16] ^ 1);
  assign comp[288] = ~(|w288);
  wire [74-1:0] w289;
  assign w289[0] = |(datain[311:308] ^ 9);
  assign w289[1] = |(datain[307:304] ^ 4);
  assign w289[2] = |(datain[303:300] ^ 4);
  assign w289[3] = |(datain[299:296] ^ 11);
  assign w289[4] = |(datain[295:292] ^ 1);
  assign w289[5] = |(datain[291:288] ^ 10);
  assign w289[6] = |(datain[287:284] ^ 12);
  assign w289[7] = |(datain[283:280] ^ 1);
  assign w289[8] = |(datain[279:276] ^ 11);
  assign w289[9] = |(datain[275:272] ^ 10);
  assign w289[10] = |(datain[271:268] ^ 7);
  assign w289[11] = |(datain[267:264] ^ 1);
  assign w289[12] = |(datain[263:260] ^ 0);
  assign w289[13] = |(datain[259:256] ^ 14);
  assign w289[14] = |(datain[255:252] ^ 8);
  assign w289[15] = |(datain[251:248] ^ 5);
  assign w289[16] = |(datain[247:244] ^ 13);
  assign w289[17] = |(datain[243:240] ^ 13);
  assign w289[18] = |(datain[239:236] ^ 8);
  assign w289[19] = |(datain[235:232] ^ 1);
  assign w289[20] = |(datain[231:228] ^ 14);
  assign w289[21] = |(datain[227:224] ^ 2);
  assign w289[22] = |(datain[223:220] ^ 0);
  assign w289[23] = |(datain[219:216] ^ 6);
  assign w289[24] = |(datain[215:212] ^ 7);
  assign w289[25] = |(datain[211:208] ^ 0);
  assign w289[26] = |(datain[207:204] ^ 11);
  assign w289[27] = |(datain[203:200] ^ 0);
  assign w289[28] = |(datain[199:196] ^ 3);
  assign w289[29] = |(datain[195:192] ^ 13);
  assign w289[30] = |(datain[191:188] ^ 12);
  assign w289[31] = |(datain[187:184] ^ 13);
  assign w289[32] = |(datain[183:180] ^ 2);
  assign w289[33] = |(datain[179:176] ^ 1);
  assign w289[34] = |(datain[175:172] ^ 14);
  assign w289[35] = |(datain[171:168] ^ 9);
  assign w289[36] = |(datain[167:164] ^ 6);
  assign w289[37] = |(datain[163:160] ^ 5);
  assign w289[38] = |(datain[159:156] ^ 0);
  assign w289[39] = |(datain[155:152] ^ 2);
  assign w289[40] = |(datain[151:148] ^ 8);
  assign w289[41] = |(datain[147:144] ^ 10);
  assign w289[42] = |(datain[143:140] ^ 14);
  assign w289[43] = |(datain[139:136] ^ 13);
  assign w289[44] = |(datain[135:132] ^ 1);
  assign w289[45] = |(datain[131:128] ^ 1);
  assign w289[46] = |(datain[127:124] ^ 8);
  assign w289[47] = |(datain[123:120] ^ 0);
  assign w289[48] = |(datain[119:116] ^ 15);
  assign w289[49] = |(datain[115:112] ^ 12);
  assign w289[50] = |(datain[111:108] ^ 3);
  assign w289[51] = |(datain[107:104] ^ 10);
  assign w289[52] = |(datain[103:100] ^ 7);
  assign w289[53] = |(datain[99:96] ^ 4);
  assign w289[54] = |(datain[95:92] ^ 0);
  assign w289[55] = |(datain[91:88] ^ 3);
  assign w289[56] = |(datain[87:84] ^ 14);
  assign w289[57] = |(datain[83:80] ^ 9);
  assign w289[58] = |(datain[79:76] ^ 0);
  assign w289[59] = |(datain[75:72] ^ 8);
  assign w289[60] = |(datain[71:68] ^ 0);
  assign w289[61] = |(datain[67:64] ^ 13);
  assign w289[62] = |(datain[63:60] ^ 3);
  assign w289[63] = |(datain[59:56] ^ 14);
  assign w289[64] = |(datain[55:52] ^ 6);
  assign w289[65] = |(datain[51:48] ^ 6);
  assign w289[66] = |(datain[47:44] ^ 8);
  assign w289[67] = |(datain[43:40] ^ 11);
  assign w289[68] = |(datain[39:36] ^ 1);
  assign w289[69] = |(datain[35:32] ^ 13);
  assign w289[70] = |(datain[31:28] ^ 14);
  assign w289[71] = |(datain[27:24] ^ 9);
  assign w289[72] = |(datain[23:20] ^ 0);
  assign w289[73] = |(datain[19:16] ^ 1);
  assign comp[289] = ~(|w289);
  wire [76-1:0] w290;
  assign w290[0] = |(datain[311:308] ^ 2);
  assign w290[1] = |(datain[307:304] ^ 1);
  assign w290[2] = |(datain[303:300] ^ 2);
  assign w290[3] = |(datain[299:296] ^ 13);
  assign w290[4] = |(datain[295:292] ^ 0);
  assign w290[5] = |(datain[291:288] ^ 3);
  assign w290[6] = |(datain[287:284] ^ 0);
  assign w290[7] = |(datain[283:280] ^ 0);
  assign w290[8] = |(datain[279:276] ^ 12);
  assign w290[9] = |(datain[275:272] ^ 6);
  assign w290[10] = |(datain[271:268] ^ 0);
  assign w290[11] = |(datain[267:264] ^ 6);
  assign w290[12] = |(datain[263:260] ^ 10);
  assign w290[13] = |(datain[259:256] ^ 14);
  assign w290[14] = |(datain[255:252] ^ 0);
  assign w290[15] = |(datain[251:248] ^ 2);
  assign w290[16] = |(datain[247:244] ^ 14);
  assign w290[17] = |(datain[243:240] ^ 9);
  assign w290[18] = |(datain[239:236] ^ 10);
  assign w290[19] = |(datain[235:232] ^ 3);
  assign w290[20] = |(datain[231:228] ^ 10);
  assign w290[21] = |(datain[227:224] ^ 15);
  assign w290[22] = |(datain[223:220] ^ 0);
  assign w290[23] = |(datain[219:216] ^ 2);
  assign w290[24] = |(datain[215:212] ^ 11);
  assign w290[25] = |(datain[211:208] ^ 4);
  assign w290[26] = |(datain[207:204] ^ 4);
  assign w290[27] = |(datain[203:200] ^ 0);
  assign w290[28] = |(datain[199:196] ^ 11);
  assign w290[29] = |(datain[195:192] ^ 9);
  assign w290[30] = |(datain[191:188] ^ 10);
  assign w290[31] = |(datain[187:184] ^ 2);
  assign w290[32] = |(datain[183:180] ^ 0);
  assign w290[33] = |(datain[179:176] ^ 2);
  assign w290[34] = |(datain[175:172] ^ 9);
  assign w290[35] = |(datain[171:168] ^ 9);
  assign w290[36] = |(datain[167:164] ^ 12);
  assign w290[37] = |(datain[163:160] ^ 13);
  assign w290[38] = |(datain[159:156] ^ 2);
  assign w290[39] = |(datain[155:152] ^ 1);
  assign w290[40] = |(datain[151:148] ^ 11);
  assign w290[41] = |(datain[147:144] ^ 8);
  assign w290[42] = |(datain[143:140] ^ 0);
  assign w290[43] = |(datain[139:136] ^ 0);
  assign w290[44] = |(datain[135:132] ^ 4);
  assign w290[45] = |(datain[131:128] ^ 2);
  assign w290[46] = |(datain[127:124] ^ 2);
  assign w290[47] = |(datain[123:120] ^ 11);
  assign w290[48] = |(datain[119:116] ^ 12);
  assign w290[49] = |(datain[115:112] ^ 9);
  assign w290[50] = |(datain[111:108] ^ 12);
  assign w290[51] = |(datain[107:104] ^ 13);
  assign w290[52] = |(datain[103:100] ^ 2);
  assign w290[53] = |(datain[99:96] ^ 1);
  assign w290[54] = |(datain[95:92] ^ 11);
  assign w290[55] = |(datain[91:88] ^ 4);
  assign w290[56] = |(datain[87:84] ^ 4);
  assign w290[57] = |(datain[83:80] ^ 0);
  assign w290[58] = |(datain[79:76] ^ 11);
  assign w290[59] = |(datain[75:72] ^ 9);
  assign w290[60] = |(datain[71:68] ^ 1);
  assign w290[61] = |(datain[67:64] ^ 10);
  assign w290[62] = |(datain[63:60] ^ 0);
  assign w290[63] = |(datain[59:56] ^ 0);
  assign w290[64] = |(datain[55:52] ^ 11);
  assign w290[65] = |(datain[51:48] ^ 10);
  assign w290[66] = |(datain[47:44] ^ 10);
  assign w290[67] = |(datain[43:40] ^ 14);
  assign w290[68] = |(datain[39:36] ^ 0);
  assign w290[69] = |(datain[35:32] ^ 2);
  assign w290[70] = |(datain[31:28] ^ 12);
  assign w290[71] = |(datain[27:24] ^ 13);
  assign w290[72] = |(datain[23:20] ^ 2);
  assign w290[73] = |(datain[19:16] ^ 1);
  assign w290[74] = |(datain[15:12] ^ 11);
  assign w290[75] = |(datain[11:8] ^ 8);
  assign comp[290] = ~(|w290);
  wire [68-1:0] w291;
  assign w291[0] = |(datain[311:308] ^ 0);
  assign w291[1] = |(datain[307:304] ^ 3);
  assign w291[2] = |(datain[303:300] ^ 10);
  assign w291[3] = |(datain[299:296] ^ 3);
  assign w291[4] = |(datain[295:292] ^ 12);
  assign w291[5] = |(datain[291:288] ^ 8);
  assign w291[6] = |(datain[287:284] ^ 0);
  assign w291[7] = |(datain[283:280] ^ 3);
  assign w291[8] = |(datain[279:276] ^ 12);
  assign w291[9] = |(datain[275:272] ^ 7);
  assign w291[10] = |(datain[271:268] ^ 0);
  assign w291[11] = |(datain[267:264] ^ 6);
  assign w291[12] = |(datain[263:260] ^ 12);
  assign w291[13] = |(datain[259:256] ^ 12);
  assign w291[14] = |(datain[255:252] ^ 0);
  assign w291[15] = |(datain[251:248] ^ 3);
  assign w291[16] = |(datain[247:244] ^ 12);
  assign w291[17] = |(datain[243:240] ^ 5);
  assign w291[18] = |(datain[239:236] ^ 8);
  assign w291[19] = |(datain[235:232] ^ 10);
  assign w291[20] = |(datain[231:228] ^ 11);
  assign w291[21] = |(datain[227:224] ^ 10);
  assign w291[22] = |(datain[223:220] ^ 0);
  assign w291[23] = |(datain[219:216] ^ 0);
  assign w291[24] = |(datain[215:212] ^ 0);
  assign w291[25] = |(datain[211:208] ^ 1);
  assign w291[26] = |(datain[207:204] ^ 11);
  assign w291[27] = |(datain[203:200] ^ 9);
  assign w291[28] = |(datain[199:196] ^ 11);
  assign w291[29] = |(datain[195:192] ^ 6);
  assign w291[30] = |(datain[191:188] ^ 0);
  assign w291[31] = |(datain[187:184] ^ 2);
  assign w291[32] = |(datain[183:180] ^ 11);
  assign w291[33] = |(datain[179:176] ^ 4);
  assign w291[34] = |(datain[175:172] ^ 4);
  assign w291[35] = |(datain[171:168] ^ 0);
  assign w291[36] = |(datain[167:164] ^ 5);
  assign w291[37] = |(datain[163:160] ^ 0);
  assign w291[38] = |(datain[159:156] ^ 12);
  assign w291[39] = |(datain[155:152] ^ 13);
  assign w291[40] = |(datain[151:148] ^ 2);
  assign w291[41] = |(datain[147:144] ^ 1);
  assign w291[42] = |(datain[143:140] ^ 14);
  assign w291[43] = |(datain[139:136] ^ 8);
  assign w291[44] = |(datain[135:132] ^ 2);
  assign w291[45] = |(datain[131:128] ^ 14);
  assign w291[46] = |(datain[127:124] ^ 15);
  assign w291[47] = |(datain[123:120] ^ 15);
  assign w291[48] = |(datain[119:116] ^ 11);
  assign w291[49] = |(datain[115:112] ^ 9);
  assign w291[50] = |(datain[111:108] ^ 0);
  assign w291[51] = |(datain[107:104] ^ 0);
  assign w291[52] = |(datain[103:100] ^ 0);
  assign w291[53] = |(datain[99:96] ^ 2);
  assign w291[54] = |(datain[95:92] ^ 15);
  assign w291[55] = |(datain[91:88] ^ 7);
  assign w291[56] = |(datain[87:84] ^ 15);
  assign w291[57] = |(datain[83:80] ^ 1);
  assign w291[58] = |(datain[79:76] ^ 8);
  assign w291[59] = |(datain[75:72] ^ 5);
  assign w291[60] = |(datain[71:68] ^ 13);
  assign w291[61] = |(datain[67:64] ^ 2);
  assign w291[62] = |(datain[63:60] ^ 7);
  assign w291[63] = |(datain[59:56] ^ 4);
  assign w291[64] = |(datain[55:52] ^ 0);
  assign w291[65] = |(datain[51:48] ^ 1);
  assign w291[66] = |(datain[47:44] ^ 4);
  assign w291[67] = |(datain[43:40] ^ 0);
  assign comp[291] = ~(|w291);
  wire [66-1:0] w292;
  assign w292[0] = |(datain[311:308] ^ 8);
  assign w292[1] = |(datain[307:304] ^ 11);
  assign w292[2] = |(datain[303:300] ^ 0);
  assign w292[3] = |(datain[299:296] ^ 14);
  assign w292[4] = |(datain[295:292] ^ 2);
  assign w292[5] = |(datain[291:288] ^ 7);
  assign w292[6] = |(datain[287:284] ^ 0);
  assign w292[7] = |(datain[283:280] ^ 1);
  assign w292[8] = |(datain[279:276] ^ 11);
  assign w292[9] = |(datain[275:272] ^ 4);
  assign w292[10] = |(datain[271:268] ^ 4);
  assign w292[11] = |(datain[267:264] ^ 14);
  assign w292[12] = |(datain[263:260] ^ 12);
  assign w292[13] = |(datain[259:256] ^ 13);
  assign w292[14] = |(datain[255:252] ^ 2);
  assign w292[15] = |(datain[251:248] ^ 1);
  assign w292[16] = |(datain[247:244] ^ 7);
  assign w292[17] = |(datain[243:240] ^ 2);
  assign w292[18] = |(datain[239:236] ^ 0);
  assign w292[19] = |(datain[235:232] ^ 15);
  assign w292[20] = |(datain[231:228] ^ 14);
  assign w292[21] = |(datain[227:224] ^ 8);
  assign w292[22] = |(datain[223:220] ^ 6);
  assign w292[23] = |(datain[219:216] ^ 11);
  assign w292[24] = |(datain[215:212] ^ 15);
  assign w292[25] = |(datain[211:208] ^ 15);
  assign w292[26] = |(datain[207:204] ^ 14);
  assign w292[27] = |(datain[203:200] ^ 8);
  assign w292[28] = |(datain[199:196] ^ 9);
  assign w292[29] = |(datain[195:192] ^ 2);
  assign w292[30] = |(datain[191:188] ^ 15);
  assign w292[31] = |(datain[187:184] ^ 15);
  assign w292[32] = |(datain[183:180] ^ 14);
  assign w292[33] = |(datain[179:176] ^ 8);
  assign w292[34] = |(datain[175:172] ^ 9);
  assign w292[35] = |(datain[171:168] ^ 11);
  assign w292[36] = |(datain[167:164] ^ 15);
  assign w292[37] = |(datain[163:160] ^ 15);
  assign w292[38] = |(datain[159:156] ^ 11);
  assign w292[39] = |(datain[155:152] ^ 4);
  assign w292[40] = |(datain[151:148] ^ 4);
  assign w292[41] = |(datain[147:144] ^ 15);
  assign w292[42] = |(datain[143:140] ^ 12);
  assign w292[43] = |(datain[139:136] ^ 13);
  assign w292[44] = |(datain[135:132] ^ 2);
  assign w292[45] = |(datain[131:128] ^ 1);
  assign w292[46] = |(datain[127:124] ^ 7);
  assign w292[47] = |(datain[123:120] ^ 5);
  assign w292[48] = |(datain[119:116] ^ 15);
  assign w292[49] = |(datain[115:112] ^ 1);
  assign w292[50] = |(datain[111:108] ^ 14);
  assign w292[51] = |(datain[107:104] ^ 8);
  assign w292[52] = |(datain[103:100] ^ 4);
  assign w292[53] = |(datain[99:96] ^ 5);
  assign w292[54] = |(datain[95:92] ^ 15);
  assign w292[55] = |(datain[91:88] ^ 15);
  assign w292[56] = |(datain[87:84] ^ 11);
  assign w292[57] = |(datain[83:80] ^ 14);
  assign w292[58] = |(datain[79:76] ^ 9);
  assign w292[59] = |(datain[75:72] ^ 9);
  assign w292[60] = |(datain[71:68] ^ 0);
  assign w292[61] = |(datain[67:64] ^ 3);
  assign w292[62] = |(datain[63:60] ^ 12);
  assign w292[63] = |(datain[59:56] ^ 13);
  assign w292[64] = |(datain[55:52] ^ 2);
  assign w292[65] = |(datain[51:48] ^ 14);
  assign comp[292] = ~(|w292);
  wire [56-1:0] w293;
  assign w293[0] = |(datain[311:308] ^ 4);
  assign w293[1] = |(datain[307:304] ^ 8);
  assign w293[2] = |(datain[303:300] ^ 0);
  assign w293[3] = |(datain[299:296] ^ 1);
  assign w293[4] = |(datain[295:292] ^ 8);
  assign w293[5] = |(datain[291:288] ^ 11);
  assign w293[6] = |(datain[287:284] ^ 9);
  assign w293[7] = |(datain[283:280] ^ 4);
  assign w293[8] = |(datain[279:276] ^ 1);
  assign w293[9] = |(datain[275:272] ^ 6);
  assign w293[10] = |(datain[271:268] ^ 0);
  assign w293[11] = |(datain[267:264] ^ 1);
  assign w293[12] = |(datain[263:260] ^ 11);
  assign w293[13] = |(datain[259:256] ^ 9);
  assign w293[14] = |(datain[255:252] ^ 11);
  assign w293[15] = |(datain[251:248] ^ 12);
  assign w293[16] = |(datain[247:244] ^ 0);
  assign w293[17] = |(datain[243:240] ^ 0);
  assign w293[18] = |(datain[239:236] ^ 8);
  assign w293[19] = |(datain[235:232] ^ 11);
  assign w293[20] = |(datain[231:228] ^ 0);
  assign w293[21] = |(datain[227:224] ^ 7);
  assign w293[22] = |(datain[223:220] ^ 3);
  assign w293[23] = |(datain[219:216] ^ 3);
  assign w293[24] = |(datain[215:212] ^ 12);
  assign w293[25] = |(datain[211:208] ^ 2);
  assign w293[26] = |(datain[207:204] ^ 8);
  assign w293[27] = |(datain[203:200] ^ 6);
  assign w293[28] = |(datain[199:196] ^ 14);
  assign w293[29] = |(datain[195:192] ^ 0);
  assign w293[30] = |(datain[191:188] ^ 3);
  assign w293[31] = |(datain[187:184] ^ 3);
  assign w293[32] = |(datain[183:180] ^ 12);
  assign w293[33] = |(datain[179:176] ^ 2);
  assign w293[34] = |(datain[175:172] ^ 8);
  assign w293[35] = |(datain[171:168] ^ 6);
  assign w293[36] = |(datain[167:164] ^ 14);
  assign w293[37] = |(datain[163:160] ^ 0);
  assign w293[38] = |(datain[159:156] ^ 8);
  assign w293[39] = |(datain[155:152] ^ 9);
  assign w293[40] = |(datain[151:148] ^ 0);
  assign w293[41] = |(datain[147:144] ^ 7);
  assign w293[42] = |(datain[143:140] ^ 8);
  assign w293[43] = |(datain[139:136] ^ 3);
  assign w293[44] = |(datain[135:132] ^ 12);
  assign w293[45] = |(datain[131:128] ^ 3);
  assign w293[46] = |(datain[127:124] ^ 0);
  assign w293[47] = |(datain[123:120] ^ 2);
  assign w293[48] = |(datain[119:116] ^ 14);
  assign w293[49] = |(datain[115:112] ^ 2);
  assign w293[50] = |(datain[111:108] ^ 14);
  assign w293[51] = |(datain[107:104] ^ 15);
  assign w293[52] = |(datain[103:100] ^ 5);
  assign w293[53] = |(datain[99:96] ^ 11);
  assign w293[54] = |(datain[95:92] ^ 12);
  assign w293[55] = |(datain[91:88] ^ 3);
  assign comp[293] = ~(|w293);
  wire [42-1:0] w294;
  assign w294[0] = |(datain[311:308] ^ 2);
  assign w294[1] = |(datain[307:304] ^ 6);
  assign w294[2] = |(datain[303:300] ^ 0);
  assign w294[3] = |(datain[299:296] ^ 1);
  assign w294[4] = |(datain[295:292] ^ 8);
  assign w294[5] = |(datain[291:288] ^ 11);
  assign w294[6] = |(datain[287:284] ^ 15);
  assign w294[7] = |(datain[283:280] ^ 14);
  assign w294[8] = |(datain[279:276] ^ 11);
  assign w294[9] = |(datain[275:272] ^ 9);
  assign w294[10] = |(datain[271:268] ^ 7);
  assign w294[11] = |(datain[267:264] ^ 4);
  assign w294[12] = |(datain[263:260] ^ 0);
  assign w294[13] = |(datain[259:256] ^ 2);
  assign w294[14] = |(datain[255:252] ^ 14);
  assign w294[15] = |(datain[251:248] ^ 8);
  assign w294[16] = |(datain[247:244] ^ 0);
  assign w294[17] = |(datain[243:240] ^ 3);
  assign w294[18] = |(datain[239:236] ^ 0);
  assign w294[19] = |(datain[235:232] ^ 0);
  assign w294[20] = |(datain[231:228] ^ 14);
  assign w294[21] = |(datain[227:224] ^ 11);
  assign w294[22] = |(datain[223:220] ^ 0);
  assign w294[23] = |(datain[219:216] ^ 11);
  assign w294[24] = |(datain[215:212] ^ 9);
  assign w294[25] = |(datain[211:208] ^ 0);
  assign w294[26] = |(datain[207:204] ^ 10);
  assign w294[27] = |(datain[203:200] ^ 12);
  assign w294[28] = |(datain[199:196] ^ 3);
  assign w294[29] = |(datain[195:192] ^ 2);
  assign w294[30] = |(datain[191:188] ^ 0);
  assign w294[31] = |(datain[187:184] ^ 6);
  assign w294[32] = |(datain[183:180] ^ 2);
  assign w294[33] = |(datain[179:176] ^ 5);
  assign w294[34] = |(datain[175:172] ^ 0);
  assign w294[35] = |(datain[171:168] ^ 1);
  assign w294[36] = |(datain[167:164] ^ 10);
  assign w294[37] = |(datain[163:160] ^ 10);
  assign w294[38] = |(datain[159:156] ^ 14);
  assign w294[39] = |(datain[155:152] ^ 2);
  assign w294[40] = |(datain[151:148] ^ 15);
  assign w294[41] = |(datain[147:144] ^ 8);
  assign comp[294] = ~(|w294);
  wire [46-1:0] w295;
  assign w295[0] = |(datain[311:308] ^ 15);
  assign w295[1] = |(datain[307:304] ^ 5);
  assign w295[2] = |(datain[303:300] ^ 11);
  assign w295[3] = |(datain[299:296] ^ 14);
  assign w295[4] = |(datain[295:292] ^ 2);
  assign w295[5] = |(datain[291:288] ^ 6);
  assign w295[6] = |(datain[287:284] ^ 0);
  assign w295[7] = |(datain[283:280] ^ 1);
  assign w295[8] = |(datain[279:276] ^ 8);
  assign w295[9] = |(datain[275:272] ^ 9);
  assign w295[10] = |(datain[271:268] ^ 15);
  assign w295[11] = |(datain[267:264] ^ 7);
  assign w295[12] = |(datain[263:260] ^ 11);
  assign w295[13] = |(datain[259:256] ^ 9);
  assign w295[14] = |(datain[255:252] ^ 7);
  assign w295[15] = |(datain[251:248] ^ 8);
  assign w295[16] = |(datain[247:244] ^ 0);
  assign w295[17] = |(datain[243:240] ^ 2);
  assign w295[18] = |(datain[239:236] ^ 14);
  assign w295[19] = |(datain[235:232] ^ 8);
  assign w295[20] = |(datain[231:228] ^ 0);
  assign w295[21] = |(datain[227:224] ^ 3);
  assign w295[22] = |(datain[223:220] ^ 0);
  assign w295[23] = |(datain[219:216] ^ 0);
  assign w295[24] = |(datain[215:212] ^ 14);
  assign w295[25] = |(datain[211:208] ^ 9);
  assign w295[26] = |(datain[207:204] ^ 0);
  assign w295[27] = |(datain[203:200] ^ 10);
  assign w295[28] = |(datain[199:196] ^ 0);
  assign w295[29] = |(datain[195:192] ^ 0);
  assign w295[30] = |(datain[191:188] ^ 10);
  assign w295[31] = |(datain[187:184] ^ 12);
  assign w295[32] = |(datain[183:180] ^ 3);
  assign w295[33] = |(datain[179:176] ^ 2);
  assign w295[34] = |(datain[175:172] ^ 0);
  assign w295[35] = |(datain[171:168] ^ 6);
  assign w295[36] = |(datain[167:164] ^ 2);
  assign w295[37] = |(datain[163:160] ^ 5);
  assign w295[38] = |(datain[159:156] ^ 0);
  assign w295[39] = |(datain[155:152] ^ 1);
  assign w295[40] = |(datain[151:148] ^ 10);
  assign w295[41] = |(datain[147:144] ^ 10);
  assign w295[42] = |(datain[143:140] ^ 14);
  assign w295[43] = |(datain[139:136] ^ 2);
  assign w295[44] = |(datain[135:132] ^ 15);
  assign w295[45] = |(datain[131:128] ^ 8);
  assign comp[295] = ~(|w295);
  wire [58-1:0] w296;
  assign w296[0] = |(datain[311:308] ^ 8);
  assign w296[1] = |(datain[307:304] ^ 0);
  assign w296[2] = |(datain[303:300] ^ 3);
  assign w296[3] = |(datain[299:296] ^ 14);
  assign w296[4] = |(datain[295:292] ^ 0);
  assign w296[5] = |(datain[291:288] ^ 4);
  assign w296[6] = |(datain[287:284] ^ 0);
  assign w296[7] = |(datain[283:280] ^ 1);
  assign w296[8] = |(datain[279:276] ^ 11);
  assign w296[9] = |(datain[275:272] ^ 11);
  assign w296[10] = |(datain[271:268] ^ 7);
  assign w296[11] = |(datain[267:264] ^ 4);
  assign w296[12] = |(datain[263:260] ^ 1);
  assign w296[13] = |(datain[259:256] ^ 6);
  assign w296[14] = |(datain[255:252] ^ 11);
  assign w296[15] = |(datain[251:248] ^ 9);
  assign w296[16] = |(datain[247:244] ^ 1);
  assign w296[17] = |(datain[243:240] ^ 10);
  assign w296[18] = |(datain[239:236] ^ 0);
  assign w296[19] = |(datain[235:232] ^ 5);
  assign w296[20] = |(datain[231:228] ^ 9);
  assign w296[21] = |(datain[227:224] ^ 0);
  assign w296[22] = |(datain[223:220] ^ 8);
  assign w296[23] = |(datain[219:216] ^ 13);
  assign w296[24] = |(datain[215:212] ^ 3);
  assign w296[25] = |(datain[211:208] ^ 14);
  assign w296[26] = |(datain[207:204] ^ 2);
  assign w296[27] = |(datain[203:200] ^ 4);
  assign w296[28] = |(datain[199:196] ^ 0);
  assign w296[29] = |(datain[195:192] ^ 1);
  assign w296[30] = |(datain[191:188] ^ 2);
  assign w296[31] = |(datain[187:184] ^ 14);
  assign w296[32] = |(datain[183:180] ^ 8);
  assign w296[33] = |(datain[179:176] ^ 11);
  assign w296[34] = |(datain[175:172] ^ 3);
  assign w296[35] = |(datain[171:168] ^ 6);
  assign w296[36] = |(datain[167:164] ^ 0);
  assign w296[37] = |(datain[163:160] ^ 2);
  assign w296[38] = |(datain[159:156] ^ 0);
  assign w296[39] = |(datain[155:152] ^ 1);
  assign w296[40] = |(datain[151:148] ^ 2);
  assign w296[41] = |(datain[147:144] ^ 14);
  assign w296[42] = |(datain[143:140] ^ 3);
  assign w296[43] = |(datain[139:136] ^ 1);
  assign w296[44] = |(datain[135:132] ^ 3);
  assign w296[45] = |(datain[131:128] ^ 13);
  assign w296[46] = |(datain[127:124] ^ 2);
  assign w296[47] = |(datain[123:120] ^ 14);
  assign w296[48] = |(datain[119:116] ^ 3);
  assign w296[49] = |(datain[115:112] ^ 1);
  assign w296[50] = |(datain[111:108] ^ 3);
  assign w296[51] = |(datain[107:104] ^ 5);
  assign w296[52] = |(datain[103:100] ^ 4);
  assign w296[53] = |(datain[99:96] ^ 7);
  assign w296[54] = |(datain[95:92] ^ 14);
  assign w296[55] = |(datain[91:88] ^ 2);
  assign w296[56] = |(datain[87:84] ^ 15);
  assign w296[57] = |(datain[83:80] ^ 7);
  assign comp[296] = ~(|w296);
  wire [48-1:0] w297;
  assign w297[0] = |(datain[311:308] ^ 11);
  assign w297[1] = |(datain[307:304] ^ 9);
  assign w297[2] = |(datain[303:300] ^ 6);
  assign w297[3] = |(datain[299:296] ^ 15);
  assign w297[4] = |(datain[295:292] ^ 0);
  assign w297[5] = |(datain[291:288] ^ 0);
  assign w297[6] = |(datain[287:284] ^ 3);
  assign w297[7] = |(datain[283:280] ^ 2);
  assign w297[8] = |(datain[279:276] ^ 12);
  assign w297[9] = |(datain[275:272] ^ 0);
  assign w297[10] = |(datain[271:268] ^ 15);
  assign w297[11] = |(datain[267:264] ^ 3);
  assign w297[12] = |(datain[263:260] ^ 10);
  assign w297[13] = |(datain[259:256] ^ 10);
  assign w297[14] = |(datain[255:252] ^ 8);
  assign w297[15] = |(datain[251:248] ^ 13);
  assign w297[16] = |(datain[247:244] ^ 9);
  assign w297[17] = |(datain[243:240] ^ 6);
  assign w297[18] = |(datain[239:236] ^ 6);
  assign w297[19] = |(datain[235:232] ^ 3);
  assign w297[20] = |(datain[231:228] ^ 15);
  assign w297[21] = |(datain[227:224] ^ 13);
  assign w297[22] = |(datain[223:220] ^ 11);
  assign w297[23] = |(datain[219:216] ^ 4);
  assign w297[24] = |(datain[215:212] ^ 4);
  assign w297[25] = |(datain[211:208] ^ 0);
  assign w297[26] = |(datain[207:204] ^ 11);
  assign w297[27] = |(datain[203:200] ^ 9);
  assign w297[28] = |(datain[199:196] ^ 1);
  assign w297[29] = |(datain[195:192] ^ 6);
  assign w297[30] = |(datain[191:188] ^ 0);
  assign w297[31] = |(datain[187:184] ^ 3);
  assign w297[32] = |(datain[183:180] ^ 12);
  assign w297[33] = |(datain[179:176] ^ 13);
  assign w297[34] = |(datain[175:172] ^ 2);
  assign w297[35] = |(datain[171:168] ^ 1);
  assign w297[36] = |(datain[167:164] ^ 7);
  assign w297[37] = |(datain[163:160] ^ 2);
  assign w297[38] = |(datain[159:156] ^ 1);
  assign w297[39] = |(datain[155:152] ^ 3);
  assign w297[40] = |(datain[151:148] ^ 5);
  assign w297[41] = |(datain[147:144] ^ 10);
  assign w297[42] = |(datain[143:140] ^ 5);
  assign w297[43] = |(datain[139:136] ^ 9);
  assign w297[44] = |(datain[135:132] ^ 8);
  assign w297[45] = |(datain[131:128] ^ 3);
  assign w297[46] = |(datain[127:124] ^ 14);
  assign w297[47] = |(datain[123:120] ^ 1);
  assign comp[297] = ~(|w297);
  wire [46-1:0] w298;
  assign w298[0] = |(datain[311:308] ^ 4);
  assign w298[1] = |(datain[307:304] ^ 0);
  assign w298[2] = |(datain[303:300] ^ 11);
  assign w298[3] = |(datain[299:296] ^ 9);
  assign w298[4] = |(datain[295:292] ^ 8);
  assign w298[5] = |(datain[291:288] ^ 4);
  assign w298[6] = |(datain[287:284] ^ 0);
  assign w298[7] = |(datain[283:280] ^ 0);
  assign w298[8] = |(datain[279:276] ^ 9);
  assign w298[9] = |(datain[275:272] ^ 0);
  assign w298[10] = |(datain[271:268] ^ 5);
  assign w298[11] = |(datain[267:264] ^ 5);
  assign w298[12] = |(datain[263:260] ^ 5);
  assign w298[13] = |(datain[259:256] ^ 10);
  assign w298[14] = |(datain[255:252] ^ 12);
  assign w298[15] = |(datain[251:248] ^ 13);
  assign w298[16] = |(datain[247:244] ^ 2);
  assign w298[17] = |(datain[243:240] ^ 1);
  assign w298[18] = |(datain[239:236] ^ 11);
  assign w298[19] = |(datain[235:232] ^ 8);
  assign w298[20] = |(datain[231:228] ^ 0);
  assign w298[21] = |(datain[227:224] ^ 0);
  assign w298[22] = |(datain[223:220] ^ 4);
  assign w298[23] = |(datain[219:216] ^ 2);
  assign w298[24] = |(datain[215:212] ^ 3);
  assign w298[25] = |(datain[211:208] ^ 3);
  assign w298[26] = |(datain[207:204] ^ 12);
  assign w298[27] = |(datain[203:200] ^ 9);
  assign w298[28] = |(datain[199:196] ^ 3);
  assign w298[29] = |(datain[195:192] ^ 3);
  assign w298[30] = |(datain[191:188] ^ 13);
  assign w298[31] = |(datain[187:184] ^ 2);
  assign w298[32] = |(datain[183:180] ^ 12);
  assign w298[33] = |(datain[179:176] ^ 13);
  assign w298[34] = |(datain[175:172] ^ 2);
  assign w298[35] = |(datain[171:168] ^ 1);
  assign w298[36] = |(datain[167:164] ^ 5);
  assign w298[37] = |(datain[163:160] ^ 14);
  assign w298[38] = |(datain[159:156] ^ 5);
  assign w298[39] = |(datain[155:152] ^ 6);
  assign w298[40] = |(datain[151:148] ^ 8);
  assign w298[41] = |(datain[147:144] ^ 11);
  assign w298[42] = |(datain[143:140] ^ 4);
  assign w298[43] = |(datain[139:136] ^ 4);
  assign w298[44] = |(datain[135:132] ^ 1);
  assign w298[45] = |(datain[131:128] ^ 10);
  assign comp[298] = ~(|w298);
  wire [44-1:0] w299;
  assign w299[0] = |(datain[311:308] ^ 11);
  assign w299[1] = |(datain[307:304] ^ 9);
  assign w299[2] = |(datain[303:300] ^ 9);
  assign w299[3] = |(datain[299:296] ^ 13);
  assign w299[4] = |(datain[295:292] ^ 0);
  assign w299[5] = |(datain[291:288] ^ 0);
  assign w299[6] = |(datain[287:284] ^ 9);
  assign w299[7] = |(datain[283:280] ^ 0);
  assign w299[8] = |(datain[279:276] ^ 5);
  assign w299[9] = |(datain[275:272] ^ 5);
  assign w299[10] = |(datain[271:268] ^ 5);
  assign w299[11] = |(datain[267:264] ^ 10);
  assign w299[12] = |(datain[263:260] ^ 12);
  assign w299[13] = |(datain[259:256] ^ 13);
  assign w299[14] = |(datain[255:252] ^ 2);
  assign w299[15] = |(datain[251:248] ^ 1);
  assign w299[16] = |(datain[247:244] ^ 11);
  assign w299[17] = |(datain[243:240] ^ 8);
  assign w299[18] = |(datain[239:236] ^ 0);
  assign w299[19] = |(datain[235:232] ^ 0);
  assign w299[20] = |(datain[231:228] ^ 4);
  assign w299[21] = |(datain[227:224] ^ 2);
  assign w299[22] = |(datain[223:220] ^ 3);
  assign w299[23] = |(datain[219:216] ^ 3);
  assign w299[24] = |(datain[215:212] ^ 12);
  assign w299[25] = |(datain[211:208] ^ 9);
  assign w299[26] = |(datain[207:204] ^ 3);
  assign w299[27] = |(datain[203:200] ^ 3);
  assign w299[28] = |(datain[199:196] ^ 13);
  assign w299[29] = |(datain[195:192] ^ 2);
  assign w299[30] = |(datain[191:188] ^ 12);
  assign w299[31] = |(datain[187:184] ^ 13);
  assign w299[32] = |(datain[183:180] ^ 2);
  assign w299[33] = |(datain[179:176] ^ 1);
  assign w299[34] = |(datain[175:172] ^ 5);
  assign w299[35] = |(datain[171:168] ^ 14);
  assign w299[36] = |(datain[167:164] ^ 5);
  assign w299[37] = |(datain[163:160] ^ 6);
  assign w299[38] = |(datain[159:156] ^ 8);
  assign w299[39] = |(datain[155:152] ^ 11);
  assign w299[40] = |(datain[151:148] ^ 4);
  assign w299[41] = |(datain[147:144] ^ 4);
  assign w299[42] = |(datain[143:140] ^ 1);
  assign w299[43] = |(datain[139:136] ^ 10);
  assign comp[299] = ~(|w299);
  wire [46-1:0] w300;
  assign w300[0] = |(datain[311:308] ^ 4);
  assign w300[1] = |(datain[307:304] ^ 0);
  assign w300[2] = |(datain[303:300] ^ 11);
  assign w300[3] = |(datain[299:296] ^ 9);
  assign w300[4] = |(datain[295:292] ^ 10);
  assign w300[5] = |(datain[291:288] ^ 13);
  assign w300[6] = |(datain[287:284] ^ 0);
  assign w300[7] = |(datain[283:280] ^ 0);
  assign w300[8] = |(datain[279:276] ^ 9);
  assign w300[9] = |(datain[275:272] ^ 0);
  assign w300[10] = |(datain[271:268] ^ 5);
  assign w300[11] = |(datain[267:264] ^ 5);
  assign w300[12] = |(datain[263:260] ^ 5);
  assign w300[13] = |(datain[259:256] ^ 10);
  assign w300[14] = |(datain[255:252] ^ 12);
  assign w300[15] = |(datain[251:248] ^ 13);
  assign w300[16] = |(datain[247:244] ^ 2);
  assign w300[17] = |(datain[243:240] ^ 1);
  assign w300[18] = |(datain[239:236] ^ 11);
  assign w300[19] = |(datain[235:232] ^ 8);
  assign w300[20] = |(datain[231:228] ^ 0);
  assign w300[21] = |(datain[227:224] ^ 0);
  assign w300[22] = |(datain[223:220] ^ 4);
  assign w300[23] = |(datain[219:216] ^ 2);
  assign w300[24] = |(datain[215:212] ^ 3);
  assign w300[25] = |(datain[211:208] ^ 3);
  assign w300[26] = |(datain[207:204] ^ 12);
  assign w300[27] = |(datain[203:200] ^ 9);
  assign w300[28] = |(datain[199:196] ^ 3);
  assign w300[29] = |(datain[195:192] ^ 3);
  assign w300[30] = |(datain[191:188] ^ 13);
  assign w300[31] = |(datain[187:184] ^ 2);
  assign w300[32] = |(datain[183:180] ^ 12);
  assign w300[33] = |(datain[179:176] ^ 13);
  assign w300[34] = |(datain[175:172] ^ 2);
  assign w300[35] = |(datain[171:168] ^ 1);
  assign w300[36] = |(datain[167:164] ^ 5);
  assign w300[37] = |(datain[163:160] ^ 14);
  assign w300[38] = |(datain[159:156] ^ 5);
  assign w300[39] = |(datain[155:152] ^ 6);
  assign w300[40] = |(datain[151:148] ^ 8);
  assign w300[41] = |(datain[147:144] ^ 11);
  assign w300[42] = |(datain[143:140] ^ 4);
  assign w300[43] = |(datain[139:136] ^ 4);
  assign w300[44] = |(datain[135:132] ^ 1);
  assign w300[45] = |(datain[131:128] ^ 10);
  assign comp[300] = ~(|w300);
  wire [74-1:0] w301;
  assign w301[0] = |(datain[311:308] ^ 8);
  assign w301[1] = |(datain[307:304] ^ 10);
  assign w301[2] = |(datain[303:300] ^ 6);
  assign w301[3] = |(datain[299:296] ^ 6);
  assign w301[4] = |(datain[295:292] ^ 0);
  assign w301[5] = |(datain[291:288] ^ 15);
  assign w301[6] = |(datain[287:284] ^ 12);
  assign w301[7] = |(datain[283:280] ^ 13);
  assign w301[8] = |(datain[279:276] ^ 2);
  assign w301[9] = |(datain[275:272] ^ 1);
  assign w301[10] = |(datain[271:268] ^ 5);
  assign w301[11] = |(datain[267:264] ^ 9);
  assign w301[12] = |(datain[263:260] ^ 5);
  assign w301[13] = |(datain[259:256] ^ 10);
  assign w301[14] = |(datain[255:252] ^ 5);
  assign w301[15] = |(datain[251:248] ^ 8);
  assign w301[16] = |(datain[247:244] ^ 3);
  assign w301[17] = |(datain[243:240] ^ 2);
  assign w301[18] = |(datain[239:236] ^ 12);
  assign w301[19] = |(datain[235:232] ^ 0);
  assign w301[20] = |(datain[231:228] ^ 12);
  assign w301[21] = |(datain[227:224] ^ 13);
  assign w301[22] = |(datain[223:220] ^ 2);
  assign w301[23] = |(datain[219:216] ^ 1);
  assign w301[24] = |(datain[215:212] ^ 8);
  assign w301[25] = |(datain[211:208] ^ 11);
  assign w301[26] = |(datain[207:204] ^ 13);
  assign w301[27] = |(datain[203:200] ^ 7);
  assign w301[28] = |(datain[199:196] ^ 11);
  assign w301[29] = |(datain[195:192] ^ 0);
  assign w301[30] = |(datain[191:188] ^ 14);
  assign w301[31] = |(datain[187:184] ^ 9);
  assign w301[32] = |(datain[183:180] ^ 10);
  assign w301[33] = |(datain[179:176] ^ 10);
  assign w301[34] = |(datain[175:172] ^ 8);
  assign w301[35] = |(datain[171:168] ^ 11);
  assign w301[36] = |(datain[167:164] ^ 4);
  assign w301[37] = |(datain[163:160] ^ 4);
  assign w301[38] = |(datain[159:156] ^ 1);
  assign w301[39] = |(datain[155:152] ^ 10);
  assign w301[40] = |(datain[151:148] ^ 2);
  assign w301[41] = |(datain[147:144] ^ 13);
  assign w301[42] = |(datain[143:140] ^ 0);
  assign w301[43] = |(datain[139:136] ^ 3);
  assign w301[44] = |(datain[135:132] ^ 0);
  assign w301[45] = |(datain[131:128] ^ 0);
  assign w301[46] = |(datain[127:124] ^ 10);
  assign w301[47] = |(datain[123:120] ^ 11);
  assign w301[48] = |(datain[119:116] ^ 11);
  assign w301[49] = |(datain[115:112] ^ 0);
  assign w301[50] = |(datain[111:108] ^ 10);
  assign w301[51] = |(datain[107:104] ^ 13);
  assign w301[52] = |(datain[103:100] ^ 10);
  assign w301[53] = |(datain[99:96] ^ 10);
  assign w301[54] = |(datain[95:92] ^ 8);
  assign w301[55] = |(datain[91:88] ^ 11);
  assign w301[56] = |(datain[87:84] ^ 15);
  assign w301[57] = |(datain[83:80] ^ 10);
  assign w301[58] = |(datain[79:76] ^ 11);
  assign w301[59] = |(datain[75:72] ^ 1);
  assign w301[60] = |(datain[71:68] ^ 0);
  assign w301[61] = |(datain[67:64] ^ 4);
  assign w301[62] = |(datain[63:60] ^ 8);
  assign w301[63] = |(datain[59:56] ^ 10);
  assign w301[64] = |(datain[55:52] ^ 6);
  assign w301[65] = |(datain[51:48] ^ 6);
  assign w301[66] = |(datain[47:44] ^ 0);
  assign w301[67] = |(datain[43:40] ^ 15);
  assign w301[68] = |(datain[39:36] ^ 12);
  assign w301[69] = |(datain[35:32] ^ 13);
  assign w301[70] = |(datain[31:28] ^ 2);
  assign w301[71] = |(datain[27:24] ^ 1);
  assign w301[72] = |(datain[23:20] ^ 14);
  assign w301[73] = |(datain[19:16] ^ 11);
  assign comp[301] = ~(|w301);
  wire [42-1:0] w302;
  assign w302[0] = |(datain[311:308] ^ 7);
  assign w302[1] = |(datain[307:304] ^ 4);
  assign w302[2] = |(datain[303:300] ^ 0);
  assign w302[3] = |(datain[299:296] ^ 15);
  assign w302[4] = |(datain[295:292] ^ 8);
  assign w302[5] = |(datain[291:288] ^ 0);
  assign w302[6] = |(datain[287:284] ^ 15);
  assign w302[7] = |(datain[283:280] ^ 12);
  assign w302[8] = |(datain[279:276] ^ 4);
  assign w302[9] = |(datain[275:272] ^ 1);
  assign w302[10] = |(datain[271:268] ^ 7);
  assign w302[11] = |(datain[267:264] ^ 4);
  assign w302[12] = |(datain[263:260] ^ 1);
  assign w302[13] = |(datain[259:256] ^ 11);
  assign w302[14] = |(datain[255:252] ^ 8);
  assign w302[15] = |(datain[251:248] ^ 0);
  assign w302[16] = |(datain[247:244] ^ 15);
  assign w302[17] = |(datain[243:240] ^ 12);
  assign w302[18] = |(datain[239:236] ^ 1);
  assign w302[19] = |(datain[235:232] ^ 3);
  assign w302[20] = |(datain[231:228] ^ 7);
  assign w302[21] = |(datain[227:224] ^ 4);
  assign w302[22] = |(datain[223:220] ^ 1);
  assign w302[23] = |(datain[219:216] ^ 6);
  assign w302[24] = |(datain[215:212] ^ 3);
  assign w302[25] = |(datain[211:208] ^ 13);
  assign w302[26] = |(datain[207:204] ^ 0);
  assign w302[27] = |(datain[203:200] ^ 0);
  assign w302[28] = |(datain[199:196] ^ 4);
  assign w302[29] = |(datain[195:192] ^ 11);
  assign w302[30] = |(datain[191:188] ^ 7);
  assign w302[31] = |(datain[187:184] ^ 4);
  assign w302[32] = |(datain[183:180] ^ 0);
  assign w302[33] = |(datain[179:176] ^ 6);
  assign w302[34] = |(datain[175:172] ^ 9);
  assign w302[35] = |(datain[171:168] ^ 13);
  assign w302[36] = |(datain[167:164] ^ 2);
  assign w302[37] = |(datain[163:160] ^ 14);
  assign w302[38] = |(datain[159:156] ^ 15);
  assign w302[39] = |(datain[155:152] ^ 15);
  assign w302[40] = |(datain[151:148] ^ 2);
  assign w302[41] = |(datain[147:144] ^ 14);
  assign comp[302] = ~(|w302);
  wire [28-1:0] w303;
  assign w303[0] = |(datain[311:308] ^ 0);
  assign w303[1] = |(datain[307:304] ^ 12);
  assign w303[2] = |(datain[303:300] ^ 11);
  assign w303[3] = |(datain[299:296] ^ 8);
  assign w303[4] = |(datain[295:292] ^ 0);
  assign w303[5] = |(datain[291:288] ^ 0);
  assign w303[6] = |(datain[287:284] ^ 4);
  assign w303[7] = |(datain[283:280] ^ 11);
  assign w303[8] = |(datain[279:276] ^ 11);
  assign w303[9] = |(datain[275:272] ^ 10);
  assign w303[10] = |(datain[271:268] ^ 11);
  assign w303[11] = |(datain[267:264] ^ 0);
  assign w303[12] = |(datain[263:260] ^ 1);
  assign w303[13] = |(datain[259:256] ^ 2);
  assign w303[14] = |(datain[255:252] ^ 12);
  assign w303[15] = |(datain[251:248] ^ 13);
  assign w303[16] = |(datain[247:244] ^ 2);
  assign w303[17] = |(datain[243:240] ^ 1);
  assign w303[18] = |(datain[239:236] ^ 11);
  assign w303[19] = |(datain[235:232] ^ 4);
  assign w303[20] = |(datain[231:228] ^ 0);
  assign w303[21] = |(datain[227:224] ^ 2);
  assign w303[22] = |(datain[223:220] ^ 11);
  assign w303[23] = |(datain[219:216] ^ 2);
  assign w303[24] = |(datain[215:212] ^ 0);
  assign w303[25] = |(datain[211:208] ^ 7);
  assign w303[26] = |(datain[207:204] ^ 12);
  assign w303[27] = |(datain[203:200] ^ 13);
  assign comp[303] = ~(|w303);
  wire [32-1:0] w304;
  assign w304[0] = |(datain[311:308] ^ 11);
  assign w304[1] = |(datain[307:304] ^ 4);
  assign w304[2] = |(datain[303:300] ^ 15);
  assign w304[3] = |(datain[299:296] ^ 15);
  assign w304[4] = |(datain[295:292] ^ 12);
  assign w304[5] = |(datain[291:288] ^ 13);
  assign w304[6] = |(datain[287:284] ^ 1);
  assign w304[7] = |(datain[283:280] ^ 3);
  assign w304[8] = |(datain[279:276] ^ 7);
  assign w304[9] = |(datain[275:272] ^ 2);
  assign w304[10] = |(datain[271:268] ^ 1);
  assign w304[11] = |(datain[267:264] ^ 8);
  assign w304[12] = |(datain[263:260] ^ 9);
  assign w304[13] = |(datain[259:256] ^ 12);
  assign w304[14] = |(datain[255:252] ^ 11);
  assign w304[15] = |(datain[251:248] ^ 15);
  assign w304[16] = |(datain[247:244] ^ 0);
  assign w304[17] = |(datain[243:240] ^ 0);
  assign w304[18] = |(datain[239:236] ^ 0);
  assign w304[19] = |(datain[235:232] ^ 1);
  assign w304[20] = |(datain[231:228] ^ 2);
  assign w304[21] = |(datain[227:224] ^ 14);
  assign w304[22] = |(datain[223:220] ^ 8);
  assign w304[23] = |(datain[219:216] ^ 11);
  assign w304[24] = |(datain[215:212] ^ 3);
  assign w304[25] = |(datain[211:208] ^ 6);
  assign w304[26] = |(datain[207:204] ^ 6);
  assign w304[27] = |(datain[203:200] ^ 2);
  assign w304[28] = |(datain[199:196] ^ 0);
  assign w304[29] = |(datain[195:192] ^ 3);
  assign w304[30] = |(datain[191:188] ^ 0);
  assign w304[31] = |(datain[187:184] ^ 3);
  assign comp[304] = ~(|w304);
  wire [76-1:0] w305;
  assign w305[0] = |(datain[311:308] ^ 0);
  assign w305[1] = |(datain[307:304] ^ 1);
  assign w305[2] = |(datain[303:300] ^ 11);
  assign w305[3] = |(datain[299:296] ^ 4);
  assign w305[4] = |(datain[295:292] ^ 4);
  assign w305[5] = |(datain[291:288] ^ 14);
  assign w305[6] = |(datain[287:284] ^ 12);
  assign w305[7] = |(datain[283:280] ^ 13);
  assign w305[8] = |(datain[279:276] ^ 2);
  assign w305[9] = |(datain[275:272] ^ 1);
  assign w305[10] = |(datain[271:268] ^ 14);
  assign w305[11] = |(datain[267:264] ^ 4);
  assign w305[12] = |(datain[263:260] ^ 4);
  assign w305[13] = |(datain[259:256] ^ 0);
  assign w305[14] = |(datain[255:252] ^ 10);
  assign w305[15] = |(datain[251:248] ^ 8);
  assign w305[16] = |(datain[247:244] ^ 0);
  assign w305[17] = |(datain[243:240] ^ 1);
  assign w305[18] = |(datain[239:236] ^ 7);
  assign w305[19] = |(datain[235:232] ^ 4);
  assign w305[20] = |(datain[231:228] ^ 1);
  assign w305[21] = |(datain[227:224] ^ 12);
  assign w305[22] = |(datain[223:220] ^ 11);
  assign w305[23] = |(datain[219:216] ^ 10);
  assign w305[24] = |(datain[215:212] ^ 9);
  assign w305[25] = |(datain[211:208] ^ 14);
  assign w305[26] = |(datain[207:204] ^ 0);
  assign w305[27] = |(datain[203:200] ^ 0);
  assign w305[28] = |(datain[199:196] ^ 11);
  assign w305[29] = |(datain[195:192] ^ 4);
  assign w305[30] = |(datain[191:188] ^ 3);
  assign w305[31] = |(datain[187:184] ^ 12);
  assign w305[32] = |(datain[183:180] ^ 11);
  assign w305[33] = |(datain[179:176] ^ 9);
  assign w305[34] = |(datain[175:172] ^ 2);
  assign w305[35] = |(datain[171:168] ^ 0);
  assign w305[36] = |(datain[167:164] ^ 0);
  assign w305[37] = |(datain[163:160] ^ 0);
  assign w305[38] = |(datain[159:156] ^ 12);
  assign w305[39] = |(datain[155:152] ^ 13);
  assign w305[40] = |(datain[151:148] ^ 2);
  assign w305[41] = |(datain[147:144] ^ 1);
  assign w305[42] = |(datain[143:140] ^ 9);
  assign w305[43] = |(datain[139:136] ^ 3);
  assign w305[44] = |(datain[135:132] ^ 7);
  assign w305[45] = |(datain[131:128] ^ 2);
  assign w305[46] = |(datain[127:124] ^ 0);
  assign w305[47] = |(datain[123:120] ^ 15);
  assign w305[48] = |(datain[119:116] ^ 11);
  assign w305[49] = |(datain[115:112] ^ 4);
  assign w305[50] = |(datain[111:108] ^ 4);
  assign w305[51] = |(datain[107:104] ^ 0);
  assign w305[52] = |(datain[103:100] ^ 11);
  assign w305[53] = |(datain[99:96] ^ 10);
  assign w305[54] = |(datain[95:92] ^ 0);
  assign w305[55] = |(datain[91:88] ^ 0);
  assign w305[56] = |(datain[87:84] ^ 0);
  assign w305[57] = |(datain[83:80] ^ 1);
  assign w305[58] = |(datain[79:76] ^ 11);
  assign w305[59] = |(datain[75:72] ^ 9);
  assign w305[60] = |(datain[71:68] ^ 2);
  assign w305[61] = |(datain[67:64] ^ 12);
  assign w305[62] = |(datain[63:60] ^ 0);
  assign w305[63] = |(datain[59:56] ^ 6);
  assign w305[64] = |(datain[55:52] ^ 9);
  assign w305[65] = |(datain[51:48] ^ 0);
  assign w305[66] = |(datain[47:44] ^ 12);
  assign w305[67] = |(datain[43:40] ^ 13);
  assign w305[68] = |(datain[39:36] ^ 2);
  assign w305[69] = |(datain[35:32] ^ 1);
  assign w305[70] = |(datain[31:28] ^ 11);
  assign w305[71] = |(datain[27:24] ^ 4);
  assign w305[72] = |(datain[23:20] ^ 3);
  assign w305[73] = |(datain[19:16] ^ 14);
  assign w305[74] = |(datain[15:12] ^ 12);
  assign w305[75] = |(datain[11:8] ^ 13);
  assign comp[305] = ~(|w305);
  wire [42-1:0] w306;
  assign w306[0] = |(datain[311:308] ^ 7);
  assign w306[1] = |(datain[307:304] ^ 4);
  assign w306[2] = |(datain[303:300] ^ 0);
  assign w306[3] = |(datain[299:296] ^ 3);
  assign w306[4] = |(datain[295:292] ^ 14);
  assign w306[5] = |(datain[291:288] ^ 9);
  assign w306[6] = |(datain[287:284] ^ 9);
  assign w306[7] = |(datain[283:280] ^ 14);
  assign w306[8] = |(datain[279:276] ^ 0);
  assign w306[9] = |(datain[275:272] ^ 0);
  assign w306[10] = |(datain[271:268] ^ 11);
  assign w306[11] = |(datain[267:264] ^ 8);
  assign w306[12] = |(datain[263:260] ^ 12);
  assign w306[13] = |(datain[259:256] ^ 4);
  assign w306[14] = |(datain[255:252] ^ 0);
  assign w306[15] = |(datain[251:248] ^ 13);
  assign w306[16] = |(datain[247:244] ^ 12);
  assign w306[17] = |(datain[243:240] ^ 13);
  assign w306[18] = |(datain[239:236] ^ 6);
  assign w306[19] = |(datain[235:232] ^ 0);
  assign w306[20] = |(datain[231:228] ^ 2);
  assign w306[21] = |(datain[227:224] ^ 14);
  assign w306[22] = |(datain[223:220] ^ 8);
  assign w306[23] = |(datain[219:216] ^ 9);
  assign w306[24] = |(datain[215:212] ^ 1);
  assign w306[25] = |(datain[211:208] ^ 14);
  assign w306[26] = |(datain[207:204] ^ 8);
  assign w306[27] = |(datain[203:200] ^ 8);
  assign w306[28] = |(datain[199:196] ^ 0);
  assign w306[29] = |(datain[195:192] ^ 1);
  assign w306[30] = |(datain[191:188] ^ 2);
  assign w306[31] = |(datain[187:184] ^ 14);
  assign w306[32] = |(datain[183:180] ^ 8);
  assign w306[33] = |(datain[179:176] ^ 12);
  assign w306[34] = |(datain[175:172] ^ 0);
  assign w306[35] = |(datain[171:168] ^ 6);
  assign w306[36] = |(datain[167:164] ^ 8);
  assign w306[37] = |(datain[163:160] ^ 10);
  assign w306[38] = |(datain[159:156] ^ 0);
  assign w306[39] = |(datain[155:152] ^ 1);
  assign w306[40] = |(datain[151:148] ^ 5);
  assign w306[41] = |(datain[147:144] ^ 2);
  assign comp[306] = ~(|w306);
  wire [42-1:0] w307;
  assign w307[0] = |(datain[311:308] ^ 7);
  assign w307[1] = |(datain[307:304] ^ 4);
  assign w307[2] = |(datain[303:300] ^ 2);
  assign w307[3] = |(datain[299:296] ^ 3);
  assign w307[4] = |(datain[295:292] ^ 8);
  assign w307[5] = |(datain[291:288] ^ 0);
  assign w307[6] = |(datain[287:284] ^ 15);
  assign w307[7] = |(datain[283:280] ^ 12);
  assign w307[8] = |(datain[279:276] ^ 4);
  assign w307[9] = |(datain[275:272] ^ 1);
  assign w307[10] = |(datain[271:268] ^ 7);
  assign w307[11] = |(datain[267:264] ^ 4);
  assign w307[12] = |(datain[263:260] ^ 0);
  assign w307[13] = |(datain[259:256] ^ 7);
  assign w307[14] = |(datain[255:252] ^ 14);
  assign w307[15] = |(datain[251:248] ^ 9);
  assign w307[16] = |(datain[247:244] ^ 3);
  assign w307[17] = |(datain[243:240] ^ 10);
  assign w307[18] = |(datain[239:236] ^ 0);
  assign w307[19] = |(datain[235:232] ^ 1);
  assign w307[20] = |(datain[231:228] ^ 5);
  assign w307[21] = |(datain[227:224] ^ 8);
  assign w307[22] = |(datain[223:220] ^ 0);
  assign w307[23] = |(datain[219:216] ^ 7);
  assign w307[24] = |(datain[215:212] ^ 14);
  assign w307[25] = |(datain[211:208] ^ 11);
  assign w307[26] = |(datain[207:204] ^ 15);
  assign w307[27] = |(datain[203:200] ^ 9);
  assign w307[28] = |(datain[199:196] ^ 0);
  assign w307[29] = |(datain[195:192] ^ 6);
  assign w307[30] = |(datain[191:188] ^ 5);
  assign w307[31] = |(datain[187:184] ^ 0);
  assign w307[32] = |(datain[183:180] ^ 3);
  assign w307[33] = |(datain[179:176] ^ 3);
  assign w307[34] = |(datain[175:172] ^ 12);
  assign w307[35] = |(datain[171:168] ^ 0);
  assign w307[36] = |(datain[167:164] ^ 8);
  assign w307[37] = |(datain[163:160] ^ 14);
  assign w307[38] = |(datain[159:156] ^ 12);
  assign w307[39] = |(datain[155:152] ^ 0);
  assign w307[40] = |(datain[151:148] ^ 2);
  assign w307[41] = |(datain[147:144] ^ 6);
  assign comp[307] = ~(|w307);
  wire [28-1:0] w308;
  assign w308[0] = |(datain[311:308] ^ 11);
  assign w308[1] = |(datain[307:304] ^ 9);
  assign w308[2] = |(datain[303:300] ^ 1);
  assign w308[3] = |(datain[299:296] ^ 14);
  assign w308[4] = |(datain[295:292] ^ 0);
  assign w308[5] = |(datain[291:288] ^ 0);
  assign w308[6] = |(datain[287:284] ^ 11);
  assign w308[7] = |(datain[283:280] ^ 10);
  assign w308[8] = |(datain[279:276] ^ 7);
  assign w308[9] = |(datain[275:272] ^ 13);
  assign w308[10] = |(datain[271:268] ^ 0);
  assign w308[11] = |(datain[267:264] ^ 4);
  assign w308[12] = |(datain[263:260] ^ 11);
  assign w308[13] = |(datain[259:256] ^ 4);
  assign w308[14] = |(datain[255:252] ^ 3);
  assign w308[15] = |(datain[251:248] ^ 15);
  assign w308[16] = |(datain[247:244] ^ 12);
  assign w308[17] = |(datain[243:240] ^ 13);
  assign w308[18] = |(datain[239:236] ^ 2);
  assign w308[19] = |(datain[235:232] ^ 1);
  assign w308[20] = |(datain[231:228] ^ 7);
  assign w308[21] = |(datain[227:224] ^ 2);
  assign w308[22] = |(datain[223:220] ^ 4);
  assign w308[23] = |(datain[219:216] ^ 6);
  assign w308[24] = |(datain[215:212] ^ 10);
  assign w308[25] = |(datain[211:208] ^ 1);
  assign w308[26] = |(datain[207:204] ^ 1);
  assign w308[27] = |(datain[203:200] ^ 2);
  assign comp[308] = ~(|w308);
  wire [28-1:0] w309;
  assign w309[0] = |(datain[311:308] ^ 15);
  assign w309[1] = |(datain[307:304] ^ 8);
  assign w309[2] = |(datain[303:300] ^ 15);
  assign w309[3] = |(datain[299:296] ^ 9);
  assign w309[4] = |(datain[295:292] ^ 11);
  assign w309[5] = |(datain[291:288] ^ 9);
  assign w309[6] = |(datain[287:284] ^ 1);
  assign w309[7] = |(datain[283:280] ^ 2);
  assign w309[8] = |(datain[279:276] ^ 11);
  assign w309[9] = |(datain[275:272] ^ 8);
  assign w309[10] = |(datain[271:268] ^ 11);
  assign w309[11] = |(datain[267:264] ^ 14);
  assign w309[12] = |(datain[263:260] ^ 1);
  assign w309[13] = |(datain[259:256] ^ 15);
  assign w309[14] = |(datain[255:252] ^ 13);
  assign w309[15] = |(datain[251:248] ^ 9);
  assign w309[16] = |(datain[247:244] ^ 3);
  assign w309[17] = |(datain[243:240] ^ 3);
  assign w309[18] = |(datain[239:236] ^ 15);
  assign w309[19] = |(datain[235:232] ^ 15);
  assign w309[20] = |(datain[231:228] ^ 15);
  assign w309[21] = |(datain[227:224] ^ 5);
  assign w309[22] = |(datain[223:220] ^ 15);
  assign w309[23] = |(datain[219:216] ^ 9);
  assign w309[24] = |(datain[215:212] ^ 15);
  assign w309[25] = |(datain[211:208] ^ 8);
  assign w309[26] = |(datain[207:204] ^ 15);
  assign w309[27] = |(datain[203:200] ^ 12);
  assign comp[309] = ~(|w309);
  wire [42-1:0] w310;
  assign w310[0] = |(datain[311:308] ^ 8);
  assign w310[1] = |(datain[307:304] ^ 13);
  assign w310[2] = |(datain[303:300] ^ 5);
  assign w310[3] = |(datain[299:296] ^ 6);
  assign w310[4] = |(datain[295:292] ^ 15);
  assign w310[5] = |(datain[291:288] ^ 13);
  assign w310[6] = |(datain[287:284] ^ 11);
  assign w310[7] = |(datain[283:280] ^ 4);
  assign w310[8] = |(datain[279:276] ^ 4);
  assign w310[9] = |(datain[275:272] ^ 0);
  assign w310[10] = |(datain[271:268] ^ 12);
  assign w310[11] = |(datain[267:264] ^ 13);
  assign w310[12] = |(datain[263:260] ^ 2);
  assign w310[13] = |(datain[259:256] ^ 1);
  assign w310[14] = |(datain[255:252] ^ 8);
  assign w310[15] = |(datain[251:248] ^ 15);
  assign w310[16] = |(datain[247:244] ^ 4);
  assign w310[17] = |(datain[243:240] ^ 5);
  assign w310[18] = |(datain[239:236] ^ 0);
  assign w310[19] = |(datain[235:232] ^ 2);
  assign w310[20] = |(datain[231:228] ^ 8);
  assign w310[21] = |(datain[227:224] ^ 15);
  assign w310[22] = |(datain[223:220] ^ 0);
  assign w310[23] = |(datain[219:216] ^ 5);
  assign w310[24] = |(datain[215:212] ^ 11);
  assign w310[25] = |(datain[211:208] ^ 8);
  assign w310[26] = |(datain[207:204] ^ 0);
  assign w310[27] = |(datain[203:200] ^ 1);
  assign w310[28] = |(datain[199:196] ^ 5);
  assign w310[29] = |(datain[195:192] ^ 7);
  assign w310[30] = |(datain[191:188] ^ 5);
  assign w310[31] = |(datain[187:184] ^ 10);
  assign w310[32] = |(datain[183:180] ^ 5);
  assign w310[33] = |(datain[179:176] ^ 9);
  assign w310[34] = |(datain[175:172] ^ 8);
  assign w310[35] = |(datain[171:168] ^ 0);
  assign w310[36] = |(datain[167:164] ^ 12);
  assign w310[37] = |(datain[163:160] ^ 9);
  assign w310[38] = |(datain[159:156] ^ 1);
  assign w310[39] = |(datain[155:152] ^ 15);
  assign w310[40] = |(datain[151:148] ^ 12);
  assign w310[41] = |(datain[147:144] ^ 13);
  assign comp[310] = ~(|w310);
  wire [54-1:0] w311;
  assign w311[0] = |(datain[311:308] ^ 0);
  assign w311[1] = |(datain[307:304] ^ 12);
  assign w311[2] = |(datain[303:300] ^ 0);
  assign w311[3] = |(datain[299:296] ^ 0);
  assign w311[4] = |(datain[295:292] ^ 11);
  assign w311[5] = |(datain[291:288] ^ 4);
  assign w311[6] = |(datain[287:284] ^ 4);
  assign w311[7] = |(datain[283:280] ^ 12);
  assign w311[8] = |(datain[279:276] ^ 11);
  assign w311[9] = |(datain[275:272] ^ 9);
  assign w311[10] = |(datain[271:268] ^ 7);
  assign w311[11] = |(datain[267:264] ^ 6);
  assign w311[12] = |(datain[263:260] ^ 0);
  assign w311[13] = |(datain[259:256] ^ 3);
  assign w311[14] = |(datain[255:252] ^ 2);
  assign w311[15] = |(datain[251:248] ^ 14);
  assign w311[16] = |(datain[247:244] ^ 8);
  assign w311[17] = |(datain[243:240] ^ 10);
  assign w311[18] = |(datain[239:236] ^ 0);
  assign w311[19] = |(datain[235:232] ^ 5);
  assign w311[20] = |(datain[231:228] ^ 8);
  assign w311[21] = |(datain[227:224] ^ 1);
  assign w311[22] = |(datain[223:220] ^ 15);
  assign w311[23] = |(datain[219:216] ^ 15);
  assign w311[24] = |(datain[215:212] ^ 2);
  assign w311[25] = |(datain[211:208] ^ 9);
  assign w311[26] = |(datain[207:204] ^ 0);
  assign w311[27] = |(datain[203:200] ^ 0);
  assign w311[28] = |(datain[199:196] ^ 7);
  assign w311[29] = |(datain[195:192] ^ 2);
  assign w311[30] = |(datain[191:188] ^ 0);
  assign w311[31] = |(datain[187:184] ^ 5);
  assign w311[32] = |(datain[183:180] ^ 3);
  assign w311[33] = |(datain[179:176] ^ 2);
  assign w311[34] = |(datain[175:172] ^ 12);
  assign w311[35] = |(datain[171:168] ^ 4);
  assign w311[36] = |(datain[167:164] ^ 2);
  assign w311[37] = |(datain[163:160] ^ 14);
  assign w311[38] = |(datain[159:156] ^ 8);
  assign w311[39] = |(datain[155:152] ^ 8);
  assign w311[40] = |(datain[151:148] ^ 0);
  assign w311[41] = |(datain[147:144] ^ 5);
  assign w311[42] = |(datain[143:140] ^ 13);
  assign w311[43] = |(datain[139:136] ^ 0);
  assign w311[44] = |(datain[135:132] ^ 12);
  assign w311[45] = |(datain[131:128] ^ 4);
  assign w311[46] = |(datain[127:124] ^ 0);
  assign w311[47] = |(datain[123:120] ^ 2);
  assign w311[48] = |(datain[119:116] ^ 14);
  assign w311[49] = |(datain[115:112] ^ 0);
  assign w311[50] = |(datain[111:108] ^ 4);
  assign w311[51] = |(datain[107:104] ^ 7);
  assign w311[52] = |(datain[103:100] ^ 14);
  assign w311[53] = |(datain[99:96] ^ 2);
  assign comp[311] = ~(|w311);
  wire [54-1:0] w312;
  assign w312[0] = |(datain[311:308] ^ 8);
  assign w312[1] = |(datain[307:304] ^ 11);
  assign w312[2] = |(datain[303:300] ^ 15);
  assign w312[3] = |(datain[299:296] ^ 12);
  assign w312[4] = |(datain[295:292] ^ 3);
  assign w312[5] = |(datain[291:288] ^ 6);
  assign w312[6] = |(datain[287:284] ^ 8);
  assign w312[7] = |(datain[283:280] ^ 11);
  assign w312[8] = |(datain[279:276] ^ 2);
  assign w312[9] = |(datain[275:272] ^ 13);
  assign w312[10] = |(datain[271:268] ^ 8);
  assign w312[11] = |(datain[267:264] ^ 1);
  assign w312[12] = |(datain[263:260] ^ 14);
  assign w312[13] = |(datain[259:256] ^ 13);
  assign w312[14] = |(datain[255:252] ^ 0);
  assign w312[15] = |(datain[251:248] ^ 3);
  assign w312[16] = |(datain[247:244] ^ 0);
  assign w312[17] = |(datain[243:240] ^ 1);
  assign w312[18] = |(datain[239:236] ^ 2);
  assign w312[19] = |(datain[235:232] ^ 14);
  assign w312[20] = |(datain[231:228] ^ 8);
  assign w312[21] = |(datain[227:224] ^ 0);
  assign w312[22] = |(datain[223:220] ^ 3);
  assign w312[23] = |(datain[219:216] ^ 14);
  assign w312[24] = |(datain[215:212] ^ 5);
  assign w312[25] = |(datain[211:208] ^ 11);
  assign w312[26] = |(datain[207:204] ^ 0);
  assign w312[27] = |(datain[203:200] ^ 1);
  assign w312[28] = |(datain[199:196] ^ 11);
  assign w312[29] = |(datain[195:192] ^ 9);
  assign w312[30] = |(datain[191:188] ^ 7);
  assign w312[31] = |(datain[187:184] ^ 4);
  assign w312[32] = |(datain[183:180] ^ 5);
  assign w312[33] = |(datain[179:176] ^ 5);
  assign w312[34] = |(datain[175:172] ^ 11);
  assign w312[35] = |(datain[171:168] ^ 9);
  assign w312[36] = |(datain[167:164] ^ 3);
  assign w312[37] = |(datain[163:160] ^ 3);
  assign w312[38] = |(datain[159:156] ^ 0);
  assign w312[39] = |(datain[155:152] ^ 4);
  assign w312[40] = |(datain[151:148] ^ 8);
  assign w312[41] = |(datain[147:144] ^ 13);
  assign w312[42] = |(datain[143:140] ^ 11);
  assign w312[43] = |(datain[139:136] ^ 14);
  assign w312[44] = |(datain[135:132] ^ 5);
  assign w312[45] = |(datain[131:128] ^ 11);
  assign w312[46] = |(datain[127:124] ^ 0);
  assign w312[47] = |(datain[123:120] ^ 1);
  assign w312[48] = |(datain[119:116] ^ 11);
  assign w312[49] = |(datain[115:112] ^ 10);
  assign w312[50] = |(datain[111:108] ^ 0);
  assign w312[51] = |(datain[107:104] ^ 1);
  assign w312[52] = |(datain[103:100] ^ 0);
  assign w312[53] = |(datain[99:96] ^ 0);
  assign comp[312] = ~(|w312);
  wire [30-1:0] w313;
  assign w313[0] = |(datain[311:308] ^ 13);
  assign w313[1] = |(datain[307:304] ^ 15);
  assign w313[2] = |(datain[303:300] ^ 8);
  assign w313[3] = |(datain[299:296] ^ 14);
  assign w313[4] = |(datain[295:292] ^ 12);
  assign w313[5] = |(datain[291:288] ^ 7);
  assign w313[6] = |(datain[287:284] ^ 8);
  assign w313[7] = |(datain[283:280] ^ 14);
  assign w313[8] = |(datain[279:276] ^ 13);
  assign w313[9] = |(datain[275:272] ^ 7);
  assign w313[10] = |(datain[271:268] ^ 8);
  assign w313[11] = |(datain[267:264] ^ 11);
  assign w313[12] = |(datain[263:260] ^ 15);
  assign w313[13] = |(datain[259:256] ^ 12);
  assign w313[14] = |(datain[255:252] ^ 11);
  assign w313[15] = |(datain[251:248] ^ 12);
  assign w313[16] = |(datain[247:244] ^ 12);
  assign w313[17] = |(datain[243:240] ^ 10);
  assign w313[18] = |(datain[239:236] ^ 0);
  assign w313[19] = |(datain[235:232] ^ 10);
  assign w313[20] = |(datain[231:228] ^ 15);
  assign w313[21] = |(datain[227:224] ^ 12);
  assign w313[22] = |(datain[223:220] ^ 14);
  assign w313[23] = |(datain[219:216] ^ 8);
  assign w313[24] = |(datain[215:212] ^ 0);
  assign w313[25] = |(datain[211:208] ^ 3);
  assign w313[26] = |(datain[207:204] ^ 0);
  assign w313[27] = |(datain[203:200] ^ 0);
  assign w313[28] = |(datain[199:196] ^ 14);
  assign w313[29] = |(datain[195:192] ^ 9);
  assign comp[313] = ~(|w313);
  wire [32-1:0] w314;
  assign w314[0] = |(datain[311:308] ^ 1);
  assign w314[1] = |(datain[307:304] ^ 4);
  assign w314[2] = |(datain[303:300] ^ 0);
  assign w314[3] = |(datain[299:296] ^ 0);
  assign w314[4] = |(datain[295:292] ^ 3);
  assign w314[5] = |(datain[291:288] ^ 1);
  assign w314[6] = |(datain[287:284] ^ 0);
  assign w314[7] = |(datain[283:280] ^ 4);
  assign w314[8] = |(datain[279:276] ^ 4);
  assign w314[9] = |(datain[275:272] ^ 6);
  assign w314[10] = |(datain[271:268] ^ 4);
  assign w314[11] = |(datain[267:264] ^ 6);
  assign w314[12] = |(datain[263:260] ^ 14);
  assign w314[13] = |(datain[259:256] ^ 2);
  assign w314[14] = |(datain[255:252] ^ 15);
  assign w314[15] = |(datain[251:248] ^ 2);
  assign w314[16] = |(datain[247:244] ^ 5);
  assign w314[17] = |(datain[243:240] ^ 14);
  assign w314[18] = |(datain[239:236] ^ 5);
  assign w314[19] = |(datain[235:232] ^ 9);
  assign w314[20] = |(datain[231:228] ^ 5);
  assign w314[21] = |(datain[227:224] ^ 8);
  assign w314[22] = |(datain[223:220] ^ 12);
  assign w314[23] = |(datain[219:216] ^ 3);
  assign w314[24] = |(datain[215:212] ^ 14);
  assign w314[25] = |(datain[211:208] ^ 8);
  assign w314[26] = |(datain[207:204] ^ 13);
  assign w314[27] = |(datain[203:200] ^ 15);
  assign w314[28] = |(datain[199:196] ^ 15);
  assign w314[29] = |(datain[195:192] ^ 15);
  assign w314[30] = |(datain[191:188] ^ 12);
  assign w314[31] = |(datain[187:184] ^ 13);
  assign comp[314] = ~(|w314);
  wire [76-1:0] w315;
  assign w315[0] = |(datain[311:308] ^ 11);
  assign w315[1] = |(datain[307:304] ^ 10);
  assign w315[2] = |(datain[303:300] ^ 0);
  assign w315[3] = |(datain[299:296] ^ 0);
  assign w315[4] = |(datain[295:292] ^ 0);
  assign w315[5] = |(datain[291:288] ^ 1);
  assign w315[6] = |(datain[287:284] ^ 11);
  assign w315[7] = |(datain[283:280] ^ 9);
  assign w315[8] = |(datain[279:276] ^ 2);
  assign w315[9] = |(datain[275:272] ^ 1);
  assign w315[10] = |(datain[271:268] ^ 0);
  assign w315[11] = |(datain[267:264] ^ 5);
  assign w315[12] = |(datain[263:260] ^ 12);
  assign w315[13] = |(datain[259:256] ^ 13);
  assign w315[14] = |(datain[255:252] ^ 2);
  assign w315[15] = |(datain[251:248] ^ 1);
  assign w315[16] = |(datain[247:244] ^ 11);
  assign w315[17] = |(datain[243:240] ^ 8);
  assign w315[18] = |(datain[239:236] ^ 0);
  assign w315[19] = |(datain[235:232] ^ 0);
  assign w315[20] = |(datain[231:228] ^ 4);
  assign w315[21] = |(datain[227:224] ^ 2);
  assign w315[22] = |(datain[223:220] ^ 3);
  assign w315[23] = |(datain[219:216] ^ 3);
  assign w315[24] = |(datain[215:212] ^ 12);
  assign w315[25] = |(datain[211:208] ^ 9);
  assign w315[26] = |(datain[207:204] ^ 3);
  assign w315[27] = |(datain[203:200] ^ 3);
  assign w315[28] = |(datain[199:196] ^ 13);
  assign w315[29] = |(datain[195:192] ^ 2);
  assign w315[30] = |(datain[191:188] ^ 12);
  assign w315[31] = |(datain[187:184] ^ 13);
  assign w315[32] = |(datain[183:180] ^ 2);
  assign w315[33] = |(datain[179:176] ^ 1);
  assign w315[34] = |(datain[175:172] ^ 11);
  assign w315[35] = |(datain[171:168] ^ 0);
  assign w315[36] = |(datain[167:164] ^ 14);
  assign w315[37] = |(datain[163:160] ^ 9);
  assign w315[38] = |(datain[159:156] ^ 10);
  assign w315[39] = |(datain[155:152] ^ 2);
  assign w315[40] = |(datain[151:148] ^ 1);
  assign w315[41] = |(datain[147:144] ^ 11);
  assign w315[42] = |(datain[143:140] ^ 0);
  assign w315[43] = |(datain[139:136] ^ 4);
  assign w315[44] = |(datain[135:132] ^ 10);
  assign w315[45] = |(datain[131:128] ^ 1);
  assign w315[46] = |(datain[127:124] ^ 1);
  assign w315[47] = |(datain[123:120] ^ 15);
  assign w315[48] = |(datain[119:116] ^ 0);
  assign w315[49] = |(datain[115:112] ^ 4);
  assign w315[50] = |(datain[111:108] ^ 2);
  assign w315[51] = |(datain[107:104] ^ 13);
  assign w315[52] = |(datain[103:100] ^ 0);
  assign w315[53] = |(datain[99:96] ^ 3);
  assign w315[54] = |(datain[95:92] ^ 0);
  assign w315[55] = |(datain[91:88] ^ 0);
  assign w315[56] = |(datain[87:84] ^ 10);
  assign w315[57] = |(datain[83:80] ^ 3);
  assign w315[58] = |(datain[79:76] ^ 1);
  assign w315[59] = |(datain[75:72] ^ 12);
  assign w315[60] = |(datain[71:68] ^ 0);
  assign w315[61] = |(datain[67:64] ^ 4);
  assign w315[62] = |(datain[63:60] ^ 11);
  assign w315[63] = |(datain[59:56] ^ 4);
  assign w315[64] = |(datain[55:52] ^ 4);
  assign w315[65] = |(datain[51:48] ^ 0);
  assign w315[66] = |(datain[47:44] ^ 11);
  assign w315[67] = |(datain[43:40] ^ 10);
  assign w315[68] = |(datain[39:36] ^ 1);
  assign w315[69] = |(datain[35:32] ^ 11);
  assign w315[70] = |(datain[31:28] ^ 0);
  assign w315[71] = |(datain[27:24] ^ 4);
  assign w315[72] = |(datain[23:20] ^ 11);
  assign w315[73] = |(datain[19:16] ^ 9);
  assign w315[74] = |(datain[15:12] ^ 0);
  assign w315[75] = |(datain[11:8] ^ 3);
  assign comp[315] = ~(|w315);
  wire [44-1:0] w316;
  assign w316[0] = |(datain[311:308] ^ 1);
  assign w316[1] = |(datain[307:304] ^ 14);
  assign w316[2] = |(datain[303:300] ^ 0);
  assign w316[3] = |(datain[299:296] ^ 5);
  assign w316[4] = |(datain[295:292] ^ 0);
  assign w316[5] = |(datain[291:288] ^ 0);
  assign w316[6] = |(datain[287:284] ^ 11);
  assign w316[7] = |(datain[283:280] ^ 5);
  assign w316[8] = |(datain[279:276] ^ 7);
  assign w316[9] = |(datain[275:272] ^ 4);
  assign w316[10] = |(datain[271:268] ^ 0);
  assign w316[11] = |(datain[267:264] ^ 3);
  assign w316[12] = |(datain[263:260] ^ 14);
  assign w316[13] = |(datain[259:256] ^ 9);
  assign w316[14] = |(datain[255:252] ^ 14);
  assign w316[15] = |(datain[251:248] ^ 3);
  assign w316[16] = |(datain[247:244] ^ 0);
  assign w316[17] = |(datain[243:240] ^ 0);
  assign w316[18] = |(datain[239:236] ^ 11);
  assign w316[19] = |(datain[235:232] ^ 8);
  assign w316[20] = |(datain[231:228] ^ 2);
  assign w316[21] = |(datain[227:224] ^ 4);
  assign w316[22] = |(datain[223:220] ^ 3);
  assign w316[23] = |(datain[219:216] ^ 5);
  assign w316[24] = |(datain[215:212] ^ 12);
  assign w316[25] = |(datain[211:208] ^ 13);
  assign w316[26] = |(datain[207:204] ^ 2);
  assign w316[27] = |(datain[203:200] ^ 1);
  assign w316[28] = |(datain[199:196] ^ 5);
  assign w316[29] = |(datain[195:192] ^ 2);
  assign w316[30] = |(datain[191:188] ^ 0);
  assign w316[31] = |(datain[187:184] ^ 14);
  assign w316[32] = |(datain[183:180] ^ 1);
  assign w316[33] = |(datain[179:176] ^ 15);
  assign w316[34] = |(datain[175:172] ^ 11);
  assign w316[35] = |(datain[171:168] ^ 10);
  assign w316[36] = |(datain[167:164] ^ 10);
  assign w316[37] = |(datain[163:160] ^ 8);
  assign w316[38] = |(datain[159:156] ^ 0);
  assign w316[39] = |(datain[155:152] ^ 0);
  assign w316[40] = |(datain[151:148] ^ 11);
  assign w316[41] = |(datain[147:144] ^ 8);
  assign w316[42] = |(datain[143:140] ^ 2);
  assign w316[43] = |(datain[139:136] ^ 4);
  assign comp[316] = ~(|w316);
  wire [28-1:0] w317;
  assign w317[0] = |(datain[311:308] ^ 12);
  assign w317[1] = |(datain[307:304] ^ 13);
  assign w317[2] = |(datain[303:300] ^ 2);
  assign w317[3] = |(datain[299:296] ^ 1);
  assign w317[4] = |(datain[295:292] ^ 11);
  assign w317[5] = |(datain[291:288] ^ 9);
  assign w317[6] = |(datain[287:284] ^ 1);
  assign w317[7] = |(datain[283:280] ^ 14);
  assign w317[8] = |(datain[279:276] ^ 15);
  assign w317[9] = |(datain[275:272] ^ 14);
  assign w317[10] = |(datain[271:268] ^ 7);
  assign w317[11] = |(datain[267:264] ^ 2);
  assign w317[12] = |(datain[263:260] ^ 2);
  assign w317[13] = |(datain[259:256] ^ 8);
  assign w317[14] = |(datain[255:252] ^ 8);
  assign w317[15] = |(datain[251:248] ^ 11);
  assign w317[16] = |(datain[247:244] ^ 13);
  assign w317[17] = |(datain[243:240] ^ 1);
  assign w317[18] = |(datain[239:236] ^ 11);
  assign w317[19] = |(datain[235:232] ^ 8);
  assign w317[20] = |(datain[231:228] ^ 0);
  assign w317[21] = |(datain[227:224] ^ 2);
  assign w317[22] = |(datain[223:220] ^ 3);
  assign w317[23] = |(datain[219:216] ^ 13);
  assign w317[24] = |(datain[215:212] ^ 12);
  assign w317[25] = |(datain[211:208] ^ 13);
  assign w317[26] = |(datain[207:204] ^ 2);
  assign w317[27] = |(datain[203:200] ^ 1);
  assign comp[317] = ~(|w317);
  wire [74-1:0] w318;
  assign w318[0] = |(datain[311:308] ^ 15);
  assign w318[1] = |(datain[307:304] ^ 15);
  assign w318[2] = |(datain[303:300] ^ 11);
  assign w318[3] = |(datain[299:296] ^ 15);
  assign w318[4] = |(datain[295:292] ^ 8);
  assign w318[5] = |(datain[291:288] ^ 5);
  assign w318[6] = |(datain[287:284] ^ 0);
  assign w318[7] = |(datain[283:280] ^ 1);
  assign w318[8] = |(datain[279:276] ^ 0);
  assign w318[9] = |(datain[275:272] ^ 14);
  assign w318[10] = |(datain[271:268] ^ 5);
  assign w318[11] = |(datain[267:264] ^ 7);
  assign w318[12] = |(datain[263:260] ^ 11);
  assign w318[13] = |(datain[259:256] ^ 8);
  assign w318[14] = |(datain[255:252] ^ 1);
  assign w318[15] = |(datain[251:248] ^ 0);
  assign w318[16] = |(datain[247:244] ^ 0);
  assign w318[17] = |(datain[243:240] ^ 0);
  assign w318[18] = |(datain[239:236] ^ 5);
  assign w318[19] = |(datain[235:232] ^ 0);
  assign w318[20] = |(datain[231:228] ^ 11);
  assign w318[21] = |(datain[227:224] ^ 15);
  assign w318[22] = |(datain[223:220] ^ 5);
  assign w318[23] = |(datain[219:216] ^ 2);
  assign w318[24] = |(datain[215:212] ^ 0);
  assign w318[25] = |(datain[211:208] ^ 0);
  assign w318[26] = |(datain[207:204] ^ 1);
  assign w318[27] = |(datain[203:200] ^ 14);
  assign w318[28] = |(datain[199:196] ^ 5);
  assign w318[29] = |(datain[195:192] ^ 7);
  assign w318[30] = |(datain[191:188] ^ 9);
  assign w318[31] = |(datain[187:184] ^ 10);
  assign w318[32] = |(datain[183:180] ^ 0);
  assign w318[33] = |(datain[179:176] ^ 0);
  assign w318[34] = |(datain[175:172] ^ 0);
  assign w318[35] = |(datain[171:168] ^ 0);
  assign w318[36] = |(datain[167:164] ^ 2);
  assign w318[37] = |(datain[163:160] ^ 3);
  assign w318[38] = |(datain[159:156] ^ 0);
  assign w318[39] = |(datain[155:152] ^ 0);
  assign w318[40] = |(datain[151:148] ^ 8);
  assign w318[41] = |(datain[147:144] ^ 3);
  assign w318[42] = |(datain[143:140] ^ 3);
  assign w318[43] = |(datain[139:136] ^ 14);
  assign w318[44] = |(datain[135:132] ^ 9);
  assign w318[45] = |(datain[131:128] ^ 2);
  assign w318[46] = |(datain[127:124] ^ 1);
  assign w318[47] = |(datain[123:120] ^ 9);
  assign w318[48] = |(datain[119:116] ^ 0);
  assign w318[49] = |(datain[115:112] ^ 0);
  assign w318[50] = |(datain[111:108] ^ 7);
  assign w318[51] = |(datain[107:104] ^ 5);
  assign w318[52] = |(datain[103:100] ^ 4);
  assign w318[53] = |(datain[99:96] ^ 15);
  assign w318[54] = |(datain[95:92] ^ 11);
  assign w318[55] = |(datain[91:88] ^ 15);
  assign w318[56] = |(datain[87:84] ^ 7);
  assign w318[57] = |(datain[83:80] ^ 0);
  assign w318[58] = |(datain[79:76] ^ 0);
  assign w318[59] = |(datain[75:72] ^ 0);
  assign w318[60] = |(datain[71:68] ^ 1);
  assign w318[61] = |(datain[67:64] ^ 14);
  assign w318[62] = |(datain[63:60] ^ 5);
  assign w318[63] = |(datain[59:56] ^ 7);
  assign w318[64] = |(datain[55:52] ^ 11);
  assign w318[65] = |(datain[51:48] ^ 15);
  assign w318[66] = |(datain[47:44] ^ 8);
  assign w318[67] = |(datain[43:40] ^ 8);
  assign w318[68] = |(datain[39:36] ^ 0);
  assign w318[69] = |(datain[35:32] ^ 1);
  assign w318[70] = |(datain[31:28] ^ 0);
  assign w318[71] = |(datain[27:24] ^ 14);
  assign w318[72] = |(datain[23:20] ^ 5);
  assign w318[73] = |(datain[19:16] ^ 7);
  assign comp[318] = ~(|w318);
  wire [76-1:0] w319;
  assign w319[0] = |(datain[311:308] ^ 3);
  assign w319[1] = |(datain[307:304] ^ 11);
  assign w319[2] = |(datain[303:300] ^ 0);
  assign w319[3] = |(datain[299:296] ^ 6);
  assign w319[4] = |(datain[295:292] ^ 0);
  assign w319[5] = |(datain[291:288] ^ 11);
  assign w319[6] = |(datain[287:284] ^ 0);
  assign w319[7] = |(datain[283:280] ^ 1);
  assign w319[8] = |(datain[279:276] ^ 7);
  assign w319[9] = |(datain[275:272] ^ 2);
  assign w319[10] = |(datain[271:268] ^ 2);
  assign w319[11] = |(datain[267:264] ^ 5);
  assign w319[12] = |(datain[263:260] ^ 11);
  assign w319[13] = |(datain[259:256] ^ 10);
  assign w319[14] = |(datain[255:252] ^ 0);
  assign w319[15] = |(datain[251:248] ^ 4);
  assign w319[16] = |(datain[247:244] ^ 0);
  assign w319[17] = |(datain[243:240] ^ 3);
  assign w319[18] = |(datain[239:236] ^ 11);
  assign w319[19] = |(datain[235:232] ^ 4);
  assign w319[20] = |(datain[231:228] ^ 4);
  assign w319[21] = |(datain[227:224] ^ 0);
  assign w319[22] = |(datain[223:220] ^ 2);
  assign w319[23] = |(datain[219:216] ^ 14);
  assign w319[24] = |(datain[215:212] ^ 8);
  assign w319[25] = |(datain[211:208] ^ 11);
  assign w319[26] = |(datain[207:204] ^ 0);
  assign w319[27] = |(datain[203:200] ^ 14);
  assign w319[28] = |(datain[199:196] ^ 0);
  assign w319[29] = |(datain[195:192] ^ 11);
  assign w319[30] = |(datain[191:188] ^ 0);
  assign w319[31] = |(datain[187:184] ^ 1);
  assign w319[32] = |(datain[183:180] ^ 12);
  assign w319[33] = |(datain[179:176] ^ 13);
  assign w319[34] = |(datain[175:172] ^ 2);
  assign w319[35] = |(datain[171:168] ^ 1);
  assign w319[36] = |(datain[167:164] ^ 7);
  assign w319[37] = |(datain[163:160] ^ 2);
  assign w319[38] = |(datain[159:156] ^ 1);
  assign w319[39] = |(datain[155:152] ^ 7);
  assign w319[40] = |(datain[151:148] ^ 11);
  assign w319[41] = |(datain[147:144] ^ 8);
  assign w319[42] = |(datain[143:140] ^ 0);
  assign w319[43] = |(datain[139:136] ^ 0);
  assign w319[44] = |(datain[135:132] ^ 4);
  assign w319[45] = |(datain[131:128] ^ 2);
  assign w319[46] = |(datain[127:124] ^ 3);
  assign w319[47] = |(datain[123:120] ^ 3);
  assign w319[48] = |(datain[119:116] ^ 12);
  assign w319[49] = |(datain[115:112] ^ 9);
  assign w319[50] = |(datain[111:108] ^ 3);
  assign w319[51] = |(datain[107:104] ^ 3);
  assign w319[52] = |(datain[103:100] ^ 13);
  assign w319[53] = |(datain[99:96] ^ 2);
  assign w319[54] = |(datain[95:92] ^ 12);
  assign w319[55] = |(datain[91:88] ^ 13);
  assign w319[56] = |(datain[87:84] ^ 2);
  assign w319[57] = |(datain[83:80] ^ 1);
  assign w319[58] = |(datain[79:76] ^ 7);
  assign w319[59] = |(datain[75:72] ^ 2);
  assign w319[60] = |(datain[71:68] ^ 0);
  assign w319[61] = |(datain[67:64] ^ 12);
  assign w319[62] = |(datain[63:60] ^ 11);
  assign w319[63] = |(datain[59:56] ^ 10);
  assign w319[64] = |(datain[55:52] ^ 0);
  assign w319[65] = |(datain[51:48] ^ 0);
  assign w319[66] = |(datain[47:44] ^ 0);
  assign w319[67] = |(datain[43:40] ^ 1);
  assign w319[68] = |(datain[39:36] ^ 11);
  assign w319[69] = |(datain[35:32] ^ 4);
  assign w319[70] = |(datain[31:28] ^ 4);
  assign w319[71] = |(datain[27:24] ^ 0);
  assign w319[72] = |(datain[23:20] ^ 2);
  assign w319[73] = |(datain[19:16] ^ 14);
  assign w319[74] = |(datain[15:12] ^ 8);
  assign w319[75] = |(datain[11:8] ^ 11);
  assign comp[319] = ~(|w319);
  wire [42-1:0] w320;
  assign w320[0] = |(datain[311:308] ^ 5);
  assign w320[1] = |(datain[307:304] ^ 10);
  assign w320[2] = |(datain[303:300] ^ 7);
  assign w320[3] = |(datain[299:296] ^ 5);
  assign w320[4] = |(datain[295:292] ^ 2);
  assign w320[5] = |(datain[291:288] ^ 4);
  assign w320[6] = |(datain[287:284] ^ 8);
  assign w320[7] = |(datain[283:280] ^ 11);
  assign w320[8] = |(datain[279:276] ^ 4);
  assign w320[9] = |(datain[275:272] ^ 4);
  assign w320[10] = |(datain[271:268] ^ 0);
  assign w320[11] = |(datain[267:264] ^ 8);
  assign w320[12] = |(datain[263:260] ^ 0);
  assign w320[13] = |(datain[259:256] ^ 3);
  assign w320[14] = |(datain[255:252] ^ 4);
  assign w320[15] = |(datain[251:248] ^ 4);
  assign w320[16] = |(datain[247:244] ^ 1);
  assign w320[17] = |(datain[243:240] ^ 6);
  assign w320[18] = |(datain[239:236] ^ 11);
  assign w320[19] = |(datain[235:232] ^ 9);
  assign w320[20] = |(datain[231:228] ^ 1);
  assign w320[21] = |(datain[227:224] ^ 0);
  assign w320[22] = |(datain[223:220] ^ 0);
  assign w320[23] = |(datain[219:216] ^ 0);
  assign w320[24] = |(datain[215:212] ^ 15);
  assign w320[25] = |(datain[211:208] ^ 7);
  assign w320[26] = |(datain[207:204] ^ 14);
  assign w320[27] = |(datain[203:200] ^ 1);
  assign w320[28] = |(datain[199:196] ^ 0);
  assign w320[29] = |(datain[195:192] ^ 3);
  assign w320[30] = |(datain[191:188] ^ 4);
  assign w320[31] = |(datain[187:184] ^ 4);
  assign w320[32] = |(datain[183:180] ^ 1);
  assign w320[33] = |(datain[179:176] ^ 4);
  assign w320[34] = |(datain[175:172] ^ 8);
  assign w320[35] = |(datain[171:168] ^ 3);
  assign w320[36] = |(datain[167:164] ^ 13);
  assign w320[37] = |(datain[163:160] ^ 2);
  assign w320[38] = |(datain[159:156] ^ 0);
  assign w320[39] = |(datain[155:152] ^ 0);
  assign w320[40] = |(datain[151:148] ^ 9);
  assign w320[41] = |(datain[147:144] ^ 2);
  assign comp[320] = ~(|w320);
  wire [46-1:0] w321;
  assign w321[0] = |(datain[311:308] ^ 7);
  assign w321[1] = |(datain[307:304] ^ 15);
  assign w321[2] = |(datain[303:300] ^ 3);
  assign w321[3] = |(datain[299:296] ^ 5);
  assign w321[4] = |(datain[295:292] ^ 12);
  assign w321[5] = |(datain[291:288] ^ 13);
  assign w321[6] = |(datain[287:284] ^ 2);
  assign w321[7] = |(datain[283:280] ^ 1);
  assign w321[8] = |(datain[279:276] ^ 8);
  assign w321[9] = |(datain[275:272] ^ 12);
  assign w321[10] = |(datain[271:268] ^ 13);
  assign w321[11] = |(datain[267:264] ^ 8);
  assign w321[12] = |(datain[263:260] ^ 8);
  assign w321[13] = |(datain[259:256] ^ 14);
  assign w321[14] = |(datain[255:252] ^ 12);
  assign w321[15] = |(datain[251:248] ^ 0);
  assign w321[16] = |(datain[247:244] ^ 8);
  assign w321[17] = |(datain[243:240] ^ 3);
  assign w321[18] = |(datain[239:236] ^ 15);
  assign w321[19] = |(datain[235:232] ^ 11);
  assign w321[20] = |(datain[231:228] ^ 15);
  assign w321[21] = |(datain[227:224] ^ 15);
  assign w321[22] = |(datain[223:220] ^ 7);
  assign w321[23] = |(datain[219:216] ^ 5);
  assign w321[24] = |(datain[215:212] ^ 0);
  assign w321[25] = |(datain[211:208] ^ 3);
  assign w321[26] = |(datain[207:204] ^ 14);
  assign w321[27] = |(datain[203:200] ^ 9);
  assign w321[28] = |(datain[199:196] ^ 9);
  assign w321[29] = |(datain[195:192] ^ 0);
  assign w321[30] = |(datain[191:188] ^ 0);
  assign w321[31] = |(datain[187:184] ^ 0);
  assign w321[32] = |(datain[183:180] ^ 11);
  assign w321[33] = |(datain[179:176] ^ 10);
  assign w321[34] = |(datain[175:172] ^ 15);
  assign w321[35] = |(datain[171:168] ^ 15);
  assign w321[36] = |(datain[167:164] ^ 15);
  assign w321[37] = |(datain[163:160] ^ 15);
  assign w321[38] = |(datain[159:156] ^ 11);
  assign w321[39] = |(datain[155:152] ^ 8);
  assign w321[40] = |(datain[151:148] ^ 7);
  assign w321[41] = |(datain[147:144] ^ 15);
  assign w321[42] = |(datain[143:140] ^ 2);
  assign w321[43] = |(datain[139:136] ^ 5);
  assign w321[44] = |(datain[135:132] ^ 12);
  assign w321[45] = |(datain[131:128] ^ 13);
  assign comp[321] = ~(|w321);
  wire [32-1:0] w322;
  assign w322[0] = |(datain[311:308] ^ 14);
  assign w322[1] = |(datain[307:304] ^ 9);
  assign w322[2] = |(datain[303:300] ^ 12);
  assign w322[3] = |(datain[299:296] ^ 12);
  assign w322[4] = |(datain[295:292] ^ 0);
  assign w322[5] = |(datain[291:288] ^ 3);
  assign w322[6] = |(datain[287:284] ^ 9);
  assign w322[7] = |(datain[283:280] ^ 0);
  assign w322[8] = |(datain[279:276] ^ 9);
  assign w322[9] = |(datain[275:272] ^ 0);
  assign w322[10] = |(datain[271:268] ^ 9);
  assign w322[11] = |(datain[267:264] ^ 0);
  assign w322[12] = |(datain[263:260] ^ 9);
  assign w322[13] = |(datain[259:256] ^ 0);
  assign w322[14] = |(datain[255:252] ^ 9);
  assign w322[15] = |(datain[251:248] ^ 0);
  assign w322[16] = |(datain[247:244] ^ 9);
  assign w322[17] = |(datain[243:240] ^ 12);
  assign w322[18] = |(datain[239:236] ^ 5);
  assign w322[19] = |(datain[235:232] ^ 0);
  assign w322[20] = |(datain[231:228] ^ 3);
  assign w322[21] = |(datain[227:224] ^ 1);
  assign w322[22] = |(datain[223:220] ^ 12);
  assign w322[23] = |(datain[219:216] ^ 0);
  assign w322[24] = |(datain[215:212] ^ 2);
  assign w322[25] = |(datain[211:208] ^ 14);
  assign w322[26] = |(datain[207:204] ^ 3);
  assign w322[27] = |(datain[203:200] ^ 8);
  assign w322[28] = |(datain[199:196] ^ 2);
  assign w322[29] = |(datain[195:192] ^ 6);
  assign w322[30] = |(datain[191:188] ^ 13);
  assign w322[31] = |(datain[187:184] ^ 10);
  assign comp[322] = ~(|w322);
  wire [30-1:0] w323;
  assign w323[0] = |(datain[311:308] ^ 2);
  assign w323[1] = |(datain[307:304] ^ 5);
  assign w323[2] = |(datain[303:300] ^ 12);
  assign w323[3] = |(datain[299:296] ^ 13);
  assign w323[4] = |(datain[295:292] ^ 2);
  assign w323[5] = |(datain[291:288] ^ 1);
  assign w323[6] = |(datain[287:284] ^ 11);
  assign w323[7] = |(datain[283:280] ^ 8);
  assign w323[8] = |(datain[279:276] ^ 2);
  assign w323[9] = |(datain[275:272] ^ 1);
  assign w323[10] = |(datain[271:268] ^ 3);
  assign w323[11] = |(datain[267:264] ^ 5);
  assign w323[12] = |(datain[263:260] ^ 12);
  assign w323[13] = |(datain[259:256] ^ 13);
  assign w323[14] = |(datain[255:252] ^ 2);
  assign w323[15] = |(datain[251:248] ^ 1);
  assign w323[16] = |(datain[247:244] ^ 8);
  assign w323[17] = |(datain[243:240] ^ 9);
  assign w323[18] = |(datain[239:236] ^ 1);
  assign w323[19] = |(datain[235:232] ^ 14);
  assign w323[20] = |(datain[231:228] ^ 14);
  assign w323[21] = |(datain[227:224] ^ 4);
  assign w323[22] = |(datain[223:220] ^ 0);
  assign w323[23] = |(datain[219:216] ^ 5);
  assign w323[24] = |(datain[215:212] ^ 8);
  assign w323[25] = |(datain[211:208] ^ 12);
  assign w323[26] = |(datain[207:204] ^ 0);
  assign w323[27] = |(datain[203:200] ^ 6);
  assign w323[28] = |(datain[199:196] ^ 14);
  assign w323[29] = |(datain[195:192] ^ 6);
  assign comp[323] = ~(|w323);
  wire [46-1:0] w324;
  assign w324[0] = |(datain[311:308] ^ 2);
  assign w324[1] = |(datain[307:304] ^ 5);
  assign w324[2] = |(datain[303:300] ^ 7);
  assign w324[3] = |(datain[299:296] ^ 5);
  assign w324[4] = |(datain[295:292] ^ 15);
  assign w324[5] = |(datain[291:288] ^ 9);
  assign w324[6] = |(datain[287:284] ^ 11);
  assign w324[7] = |(datain[283:280] ^ 10);
  assign w324[8] = |(datain[279:276] ^ 0);
  assign w324[9] = |(datain[275:272] ^ 0);
  assign w324[10] = |(datain[271:268] ^ 4);
  assign w324[11] = |(datain[267:264] ^ 2);
  assign w324[12] = |(datain[263:260] ^ 2);
  assign w324[13] = |(datain[259:256] ^ 6);
  assign w324[14] = |(datain[255:252] ^ 3);
  assign w324[15] = |(datain[251:248] ^ 11);
  assign w324[16] = |(datain[247:244] ^ 5);
  assign w324[17] = |(datain[243:240] ^ 5);
  assign w324[18] = |(datain[239:236] ^ 0);
  assign w324[19] = |(datain[235:232] ^ 1);
  assign w324[20] = |(datain[231:228] ^ 7);
  assign w324[21] = |(datain[227:224] ^ 5);
  assign w324[22] = |(datain[223:220] ^ 15);
  assign w324[23] = |(datain[219:216] ^ 0);
  assign w324[24] = |(datain[215:212] ^ 11);
  assign w324[25] = |(datain[211:208] ^ 6);
  assign w324[26] = |(datain[207:204] ^ 11);
  assign w324[27] = |(datain[203:200] ^ 10);
  assign w324[28] = |(datain[199:196] ^ 2);
  assign w324[29] = |(datain[195:192] ^ 6);
  assign w324[30] = |(datain[191:188] ^ 3);
  assign w324[31] = |(datain[187:184] ^ 10);
  assign w324[32] = |(datain[183:180] ^ 7);
  assign w324[33] = |(datain[179:176] ^ 5);
  assign w324[34] = |(datain[175:172] ^ 15);
  assign w324[35] = |(datain[171:168] ^ 11);
  assign w324[36] = |(datain[167:164] ^ 7);
  assign w324[37] = |(datain[163:160] ^ 5);
  assign w324[38] = |(datain[159:156] ^ 14);
  assign w324[39] = |(datain[155:152] ^ 8);
  assign w324[40] = |(datain[151:148] ^ 8);
  assign w324[41] = |(datain[147:144] ^ 3);
  assign w324[42] = |(datain[143:140] ^ 15);
  assign w324[43] = |(datain[139:136] ^ 9);
  assign w324[44] = |(datain[135:132] ^ 0);
  assign w324[45] = |(datain[131:128] ^ 0);
  assign comp[324] = ~(|w324);
  wire [32-1:0] w325;
  assign w325[0] = |(datain[311:308] ^ 14);
  assign w325[1] = |(datain[307:304] ^ 14);
  assign w325[2] = |(datain[303:300] ^ 11);
  assign w325[3] = |(datain[299:296] ^ 10);
  assign w325[4] = |(datain[295:292] ^ 7);
  assign w325[5] = |(datain[291:288] ^ 1);
  assign w325[6] = |(datain[287:284] ^ 0);
  assign w325[7] = |(datain[283:280] ^ 0);
  assign w325[8] = |(datain[279:276] ^ 14);
  assign w325[9] = |(datain[275:272] ^ 12);
  assign w325[10] = |(datain[271:268] ^ 3);
  assign w325[11] = |(datain[267:264] ^ 12);
  assign w325[12] = |(datain[263:260] ^ 15);
  assign w325[13] = |(datain[259:256] ^ 0);
  assign w325[14] = |(datain[255:252] ^ 7);
  assign w325[15] = |(datain[251:248] ^ 6);
  assign w325[16] = |(datain[247:244] ^ 0);
  assign w325[17] = |(datain[243:240] ^ 3);
  assign w325[18] = |(datain[239:236] ^ 14);
  assign w325[19] = |(datain[235:232] ^ 9);
  assign w325[20] = |(datain[231:228] ^ 9);
  assign w325[21] = |(datain[227:224] ^ 10);
  assign w325[22] = |(datain[223:220] ^ 0);
  assign w325[23] = |(datain[219:216] ^ 0);
  assign w325[24] = |(datain[215:212] ^ 11);
  assign w325[25] = |(datain[211:208] ^ 8);
  assign w325[26] = |(datain[207:204] ^ 7);
  assign w325[27] = |(datain[203:200] ^ 15);
  assign w325[28] = |(datain[199:196] ^ 3);
  assign w325[29] = |(datain[195:192] ^ 5);
  assign w325[30] = |(datain[191:188] ^ 12);
  assign w325[31] = |(datain[187:184] ^ 13);
  assign comp[325] = ~(|w325);
  wire [30-1:0] w326;
  assign w326[0] = |(datain[311:308] ^ 2);
  assign w326[1] = |(datain[307:304] ^ 9);
  assign w326[2] = |(datain[303:300] ^ 4);
  assign w326[3] = |(datain[299:296] ^ 13);
  assign w326[4] = |(datain[295:292] ^ 0);
  assign w326[5] = |(datain[291:288] ^ 3);
  assign w326[6] = |(datain[287:284] ^ 8);
  assign w326[7] = |(datain[283:280] ^ 9);
  assign w326[8] = |(datain[279:276] ^ 5);
  assign w326[9] = |(datain[275:272] ^ 5);
  assign w326[10] = |(datain[271:268] ^ 0);
  assign w326[11] = |(datain[267:264] ^ 2);
  assign w326[12] = |(datain[263:260] ^ 8);
  assign w326[13] = |(datain[259:256] ^ 14);
  assign w326[14] = |(datain[255:252] ^ 12);
  assign w326[15] = |(datain[251:248] ^ 2);
  assign w326[16] = |(datain[247:244] ^ 8);
  assign w326[17] = |(datain[243:240] ^ 13);
  assign w326[18] = |(datain[239:236] ^ 7);
  assign w326[19] = |(datain[235:232] ^ 7);
  assign w326[20] = |(datain[231:228] ^ 15);
  assign w326[21] = |(datain[227:224] ^ 13);
  assign w326[22] = |(datain[223:220] ^ 11);
  assign w326[23] = |(datain[219:216] ^ 9);
  assign w326[24] = |(datain[215:212] ^ 9);
  assign w326[25] = |(datain[211:208] ^ 5);
  assign w326[26] = |(datain[207:204] ^ 0);
  assign w326[27] = |(datain[203:200] ^ 4);
  assign w326[28] = |(datain[199:196] ^ 15);
  assign w326[29] = |(datain[195:192] ^ 3);
  assign comp[326] = ~(|w326);
  wire [46-1:0] w327;
  assign w327[0] = |(datain[311:308] ^ 8);
  assign w327[1] = |(datain[307:304] ^ 6);
  assign w327[2] = |(datain[303:300] ^ 3);
  assign w327[3] = |(datain[299:296] ^ 11);
  assign w327[4] = |(datain[295:292] ^ 0);
  assign w327[5] = |(datain[291:288] ^ 2);
  assign w327[6] = |(datain[287:284] ^ 11);
  assign w327[7] = |(datain[283:280] ^ 4);
  assign w327[8] = |(datain[279:276] ^ 4);
  assign w327[9] = |(datain[275:272] ^ 0);
  assign w327[10] = |(datain[271:268] ^ 11);
  assign w327[11] = |(datain[267:264] ^ 9);
  assign w327[12] = |(datain[263:260] ^ 5);
  assign w327[13] = |(datain[259:256] ^ 1);
  assign w327[14] = |(datain[255:252] ^ 0);
  assign w327[15] = |(datain[251:248] ^ 1);
  assign w327[16] = |(datain[247:244] ^ 8);
  assign w327[17] = |(datain[243:240] ^ 13);
  assign w327[18] = |(datain[239:236] ^ 9);
  assign w327[19] = |(datain[235:232] ^ 6);
  assign w327[20] = |(datain[231:228] ^ 0);
  assign w327[21] = |(datain[227:224] ^ 0);
  assign w327[22] = |(datain[223:220] ^ 0);
  assign w327[23] = |(datain[219:216] ^ 1);
  assign w327[24] = |(datain[215:212] ^ 12);
  assign w327[25] = |(datain[211:208] ^ 13);
  assign w327[26] = |(datain[207:204] ^ 2);
  assign w327[27] = |(datain[203:200] ^ 1);
  assign w327[28] = |(datain[199:196] ^ 11);
  assign w327[29] = |(datain[195:192] ^ 8);
  assign w327[30] = |(datain[191:188] ^ 0);
  assign w327[31] = |(datain[187:184] ^ 0);
  assign w327[32] = |(datain[183:180] ^ 4);
  assign w327[33] = |(datain[179:176] ^ 2);
  assign w327[34] = |(datain[175:172] ^ 3);
  assign w327[35] = |(datain[171:168] ^ 3);
  assign w327[36] = |(datain[167:164] ^ 12);
  assign w327[37] = |(datain[163:160] ^ 9);
  assign w327[38] = |(datain[159:156] ^ 3);
  assign w327[39] = |(datain[155:152] ^ 3);
  assign w327[40] = |(datain[151:148] ^ 13);
  assign w327[41] = |(datain[147:144] ^ 2);
  assign w327[42] = |(datain[143:140] ^ 12);
  assign w327[43] = |(datain[139:136] ^ 13);
  assign w327[44] = |(datain[135:132] ^ 2);
  assign w327[45] = |(datain[131:128] ^ 1);
  assign comp[327] = ~(|w327);
  wire [42-1:0] w328;
  assign w328[0] = |(datain[311:308] ^ 0);
  assign w328[1] = |(datain[307:304] ^ 2);
  assign w328[2] = |(datain[303:300] ^ 11);
  assign w328[3] = |(datain[299:296] ^ 4);
  assign w328[4] = |(datain[295:292] ^ 4);
  assign w328[5] = |(datain[291:288] ^ 0);
  assign w328[6] = |(datain[287:284] ^ 11);
  assign w328[7] = |(datain[283:280] ^ 9);
  assign w328[8] = |(datain[279:276] ^ 7);
  assign w328[9] = |(datain[275:272] ^ 11);
  assign w328[10] = |(datain[271:268] ^ 0);
  assign w328[11] = |(datain[267:264] ^ 1);
  assign w328[12] = |(datain[263:260] ^ 8);
  assign w328[13] = |(datain[259:256] ^ 13);
  assign w328[14] = |(datain[255:252] ^ 9);
  assign w328[15] = |(datain[251:248] ^ 6);
  assign w328[16] = |(datain[247:244] ^ 0);
  assign w328[17] = |(datain[243:240] ^ 0);
  assign w328[18] = |(datain[239:236] ^ 0);
  assign w328[19] = |(datain[235:232] ^ 1);
  assign w328[20] = |(datain[231:228] ^ 12);
  assign w328[21] = |(datain[227:224] ^ 13);
  assign w328[22] = |(datain[223:220] ^ 2);
  assign w328[23] = |(datain[219:216] ^ 1);
  assign w328[24] = |(datain[215:212] ^ 11);
  assign w328[25] = |(datain[211:208] ^ 8);
  assign w328[26] = |(datain[207:204] ^ 0);
  assign w328[27] = |(datain[203:200] ^ 0);
  assign w328[28] = |(datain[199:196] ^ 4);
  assign w328[29] = |(datain[195:192] ^ 2);
  assign w328[30] = |(datain[191:188] ^ 3);
  assign w328[31] = |(datain[187:184] ^ 3);
  assign w328[32] = |(datain[183:180] ^ 12);
  assign w328[33] = |(datain[179:176] ^ 9);
  assign w328[34] = |(datain[175:172] ^ 3);
  assign w328[35] = |(datain[171:168] ^ 3);
  assign w328[36] = |(datain[167:164] ^ 13);
  assign w328[37] = |(datain[163:160] ^ 2);
  assign w328[38] = |(datain[159:156] ^ 12);
  assign w328[39] = |(datain[155:152] ^ 13);
  assign w328[40] = |(datain[151:148] ^ 2);
  assign w328[41] = |(datain[147:144] ^ 1);
  assign comp[328] = ~(|w328);
  wire [74-1:0] w329;
  assign w329[0] = |(datain[311:308] ^ 0);
  assign w329[1] = |(datain[307:304] ^ 3);
  assign w329[2] = |(datain[303:300] ^ 0);
  assign w329[3] = |(datain[299:296] ^ 0);
  assign w329[4] = |(datain[295:292] ^ 8);
  assign w329[5] = |(datain[291:288] ^ 9);
  assign w329[6] = |(datain[287:284] ^ 8);
  assign w329[7] = |(datain[283:280] ^ 6);
  assign w329[8] = |(datain[279:276] ^ 2);
  assign w329[9] = |(datain[275:272] ^ 12);
  assign w329[10] = |(datain[271:268] ^ 0);
  assign w329[11] = |(datain[267:264] ^ 2);
  assign w329[12] = |(datain[263:260] ^ 11);
  assign w329[13] = |(datain[259:256] ^ 4);
  assign w329[14] = |(datain[255:252] ^ 4);
  assign w329[15] = |(datain[251:248] ^ 0);
  assign w329[16] = |(datain[247:244] ^ 11);
  assign w329[17] = |(datain[243:240] ^ 9);
  assign w329[18] = |(datain[239:236] ^ 7);
  assign w329[19] = |(datain[235:232] ^ 15);
  assign w329[20] = |(datain[231:228] ^ 0);
  assign w329[21] = |(datain[227:224] ^ 1);
  assign w329[22] = |(datain[223:220] ^ 8);
  assign w329[23] = |(datain[219:216] ^ 13);
  assign w329[24] = |(datain[215:212] ^ 9);
  assign w329[25] = |(datain[211:208] ^ 6);
  assign w329[26] = |(datain[207:204] ^ 0);
  assign w329[27] = |(datain[203:200] ^ 0);
  assign w329[28] = |(datain[199:196] ^ 0);
  assign w329[29] = |(datain[195:192] ^ 1);
  assign w329[30] = |(datain[191:188] ^ 12);
  assign w329[31] = |(datain[187:184] ^ 13);
  assign w329[32] = |(datain[183:180] ^ 2);
  assign w329[33] = |(datain[179:176] ^ 1);
  assign w329[34] = |(datain[175:172] ^ 11);
  assign w329[35] = |(datain[171:168] ^ 8);
  assign w329[36] = |(datain[167:164] ^ 0);
  assign w329[37] = |(datain[163:160] ^ 0);
  assign w329[38] = |(datain[159:156] ^ 4);
  assign w329[39] = |(datain[155:152] ^ 2);
  assign w329[40] = |(datain[151:148] ^ 3);
  assign w329[41] = |(datain[147:144] ^ 3);
  assign w329[42] = |(datain[143:140] ^ 12);
  assign w329[43] = |(datain[139:136] ^ 9);
  assign w329[44] = |(datain[135:132] ^ 3);
  assign w329[45] = |(datain[131:128] ^ 3);
  assign w329[46] = |(datain[127:124] ^ 13);
  assign w329[47] = |(datain[123:120] ^ 2);
  assign w329[48] = |(datain[119:116] ^ 12);
  assign w329[49] = |(datain[115:112] ^ 13);
  assign w329[50] = |(datain[111:108] ^ 2);
  assign w329[51] = |(datain[107:104] ^ 1);
  assign w329[52] = |(datain[103:100] ^ 11);
  assign w329[53] = |(datain[99:96] ^ 4);
  assign w329[54] = |(datain[95:92] ^ 4);
  assign w329[55] = |(datain[91:88] ^ 0);
  assign w329[56] = |(datain[87:84] ^ 11);
  assign w329[57] = |(datain[83:80] ^ 9);
  assign w329[58] = |(datain[79:76] ^ 0);
  assign w329[59] = |(datain[75:72] ^ 4);
  assign w329[60] = |(datain[71:68] ^ 0);
  assign w329[61] = |(datain[67:64] ^ 0);
  assign w329[62] = |(datain[63:60] ^ 8);
  assign w329[63] = |(datain[59:56] ^ 13);
  assign w329[64] = |(datain[55:52] ^ 9);
  assign w329[65] = |(datain[51:48] ^ 6);
  assign w329[66] = |(datain[47:44] ^ 2);
  assign w329[67] = |(datain[43:40] ^ 11);
  assign w329[68] = |(datain[39:36] ^ 0);
  assign w329[69] = |(datain[35:32] ^ 2);
  assign w329[70] = |(datain[31:28] ^ 12);
  assign w329[71] = |(datain[27:24] ^ 13);
  assign w329[72] = |(datain[23:20] ^ 2);
  assign w329[73] = |(datain[19:16] ^ 1);
  assign comp[329] = ~(|w329);
  wire [42-1:0] w330;
  assign w330[0] = |(datain[311:308] ^ 0);
  assign w330[1] = |(datain[307:304] ^ 2);
  assign w330[2] = |(datain[303:300] ^ 11);
  assign w330[3] = |(datain[299:296] ^ 4);
  assign w330[4] = |(datain[295:292] ^ 4);
  assign w330[5] = |(datain[291:288] ^ 0);
  assign w330[6] = |(datain[287:284] ^ 11);
  assign w330[7] = |(datain[283:280] ^ 9);
  assign w330[8] = |(datain[279:276] ^ 8);
  assign w330[9] = |(datain[275:272] ^ 1);
  assign w330[10] = |(datain[271:268] ^ 0);
  assign w330[11] = |(datain[267:264] ^ 1);
  assign w330[12] = |(datain[263:260] ^ 8);
  assign w330[13] = |(datain[259:256] ^ 13);
  assign w330[14] = |(datain[255:252] ^ 9);
  assign w330[15] = |(datain[251:248] ^ 6);
  assign w330[16] = |(datain[247:244] ^ 0);
  assign w330[17] = |(datain[243:240] ^ 0);
  assign w330[18] = |(datain[239:236] ^ 0);
  assign w330[19] = |(datain[235:232] ^ 1);
  assign w330[20] = |(datain[231:228] ^ 12);
  assign w330[21] = |(datain[227:224] ^ 13);
  assign w330[22] = |(datain[223:220] ^ 2);
  assign w330[23] = |(datain[219:216] ^ 1);
  assign w330[24] = |(datain[215:212] ^ 11);
  assign w330[25] = |(datain[211:208] ^ 8);
  assign w330[26] = |(datain[207:204] ^ 0);
  assign w330[27] = |(datain[203:200] ^ 0);
  assign w330[28] = |(datain[199:196] ^ 4);
  assign w330[29] = |(datain[195:192] ^ 2);
  assign w330[30] = |(datain[191:188] ^ 3);
  assign w330[31] = |(datain[187:184] ^ 3);
  assign w330[32] = |(datain[183:180] ^ 12);
  assign w330[33] = |(datain[179:176] ^ 9);
  assign w330[34] = |(datain[175:172] ^ 3);
  assign w330[35] = |(datain[171:168] ^ 3);
  assign w330[36] = |(datain[167:164] ^ 13);
  assign w330[37] = |(datain[163:160] ^ 2);
  assign w330[38] = |(datain[159:156] ^ 12);
  assign w330[39] = |(datain[155:152] ^ 13);
  assign w330[40] = |(datain[151:148] ^ 2);
  assign w330[41] = |(datain[147:144] ^ 1);
  assign comp[330] = ~(|w330);
  wire [42-1:0] w331;
  assign w331[0] = |(datain[311:308] ^ 0);
  assign w331[1] = |(datain[307:304] ^ 2);
  assign w331[2] = |(datain[303:300] ^ 8);
  assign w331[3] = |(datain[299:296] ^ 13);
  assign w331[4] = |(datain[295:292] ^ 11);
  assign w331[5] = |(datain[291:288] ^ 6);
  assign w331[6] = |(datain[287:284] ^ 0);
  assign w331[7] = |(datain[283:280] ^ 15);
  assign w331[8] = |(datain[279:276] ^ 0);
  assign w331[9] = |(datain[275:272] ^ 1);
  assign w331[10] = |(datain[271:268] ^ 14);
  assign w331[11] = |(datain[267:264] ^ 11);
  assign w331[12] = |(datain[263:260] ^ 0);
  assign w331[13] = |(datain[259:256] ^ 7);
  assign w331[14] = |(datain[255:252] ^ 10);
  assign w331[15] = |(datain[251:248] ^ 13);
  assign w331[16] = |(datain[247:244] ^ 3);
  assign w331[17] = |(datain[243:240] ^ 3);
  assign w331[18] = |(datain[239:236] ^ 12);
  assign w331[19] = |(datain[235:232] ^ 2);
  assign w331[20] = |(datain[231:228] ^ 10);
  assign w331[21] = |(datain[227:224] ^ 11);
  assign w331[22] = |(datain[223:220] ^ 14);
  assign w331[23] = |(datain[219:216] ^ 2);
  assign w331[24] = |(datain[215:212] ^ 15);
  assign w331[25] = |(datain[211:208] ^ 10);
  assign w331[26] = |(datain[207:204] ^ 12);
  assign w331[27] = |(datain[203:200] ^ 3);
  assign w331[28] = |(datain[199:196] ^ 11);
  assign w331[29] = |(datain[195:192] ^ 9);
  assign w331[30] = |(datain[191:188] ^ 8);
  assign w331[31] = |(datain[187:184] ^ 11);
  assign w331[32] = |(datain[183:180] ^ 0);
  assign w331[33] = |(datain[179:176] ^ 0);
  assign w331[34] = |(datain[175:172] ^ 8);
  assign w331[35] = |(datain[171:168] ^ 11);
  assign w331[36] = |(datain[167:164] ^ 15);
  assign w331[37] = |(datain[163:160] ^ 14);
  assign w331[38] = |(datain[159:156] ^ 14);
  assign w331[39] = |(datain[155:152] ^ 11);
  assign w331[40] = |(datain[151:148] ^ 15);
  assign w331[41] = |(datain[147:144] ^ 2);
  assign comp[331] = ~(|w331);
  wire [46-1:0] w332;
  assign w332[0] = |(datain[311:308] ^ 7);
  assign w332[1] = |(datain[307:304] ^ 11);
  assign w332[2] = |(datain[303:300] ^ 0);
  assign w332[3] = |(datain[299:296] ^ 6);
  assign w332[4] = |(datain[295:292] ^ 2);
  assign w332[5] = |(datain[291:288] ^ 14);
  assign w332[6] = |(datain[287:284] ^ 8);
  assign w332[7] = |(datain[283:280] ^ 11);
  assign w332[8] = |(datain[279:276] ^ 9);
  assign w332[9] = |(datain[275:272] ^ 12);
  assign w332[10] = |(datain[271:268] ^ 5);
  assign w332[11] = |(datain[267:264] ^ 14);
  assign w332[12] = |(datain[263:260] ^ 0);
  assign w332[13] = |(datain[259:256] ^ 7);
  assign w332[14] = |(datain[255:252] ^ 11);
  assign w332[15] = |(datain[251:248] ^ 4);
  assign w332[16] = |(datain[247:244] ^ 4);
  assign w332[17] = |(datain[243:240] ^ 0);
  assign w332[18] = |(datain[239:236] ^ 12);
  assign w332[19] = |(datain[235:232] ^ 13);
  assign w332[20] = |(datain[231:228] ^ 2);
  assign w332[21] = |(datain[227:224] ^ 1);
  assign w332[22] = |(datain[223:220] ^ 14);
  assign w332[23] = |(datain[219:216] ^ 8);
  assign w332[24] = |(datain[215:212] ^ 10);
  assign w332[25] = |(datain[211:208] ^ 15);
  assign w332[26] = |(datain[207:204] ^ 15);
  assign w332[27] = |(datain[203:200] ^ 11);
  assign w332[28] = |(datain[199:196] ^ 2);
  assign w332[29] = |(datain[195:192] ^ 14);
  assign w332[30] = |(datain[191:188] ^ 8);
  assign w332[31] = |(datain[187:184] ^ 15);
  assign w332[32] = |(datain[183:180] ^ 8);
  assign w332[33] = |(datain[179:176] ^ 4);
  assign w332[34] = |(datain[175:172] ^ 7);
  assign w332[35] = |(datain[171:168] ^ 6);
  assign w332[36] = |(datain[167:164] ^ 0);
  assign w332[37] = |(datain[163:160] ^ 7);
  assign w332[38] = |(datain[159:156] ^ 2);
  assign w332[39] = |(datain[155:152] ^ 14);
  assign w332[40] = |(datain[151:148] ^ 8);
  assign w332[41] = |(datain[147:144] ^ 15);
  assign w332[42] = |(datain[143:140] ^ 8);
  assign w332[43] = |(datain[139:136] ^ 4);
  assign w332[44] = |(datain[135:132] ^ 6);
  assign w332[45] = |(datain[131:128] ^ 13);
  assign comp[332] = ~(|w332);
  wire [28-1:0] w333;
  assign w333[0] = |(datain[311:308] ^ 10);
  assign w333[1] = |(datain[307:304] ^ 14);
  assign w333[2] = |(datain[303:300] ^ 4);
  assign w333[3] = |(datain[299:296] ^ 2);
  assign w333[4] = |(datain[295:292] ^ 6);
  assign w333[5] = |(datain[291:288] ^ 14);
  assign w333[6] = |(datain[287:284] ^ 4);
  assign w333[7] = |(datain[283:280] ^ 12);
  assign w333[8] = |(datain[279:276] ^ 7);
  assign w333[9] = |(datain[275:272] ^ 2);
  assign w333[10] = |(datain[271:268] ^ 0);
  assign w333[11] = |(datain[267:264] ^ 3);
  assign w333[12] = |(datain[263:260] ^ 4);
  assign w333[13] = |(datain[259:256] ^ 6);
  assign w333[14] = |(datain[255:252] ^ 0);
  assign w333[15] = |(datain[251:248] ^ 0);
  assign w333[16] = |(datain[247:244] ^ 0);
  assign w333[17] = |(datain[243:240] ^ 0);
  assign w333[18] = |(datain[239:236] ^ 0);
  assign w333[19] = |(datain[235:232] ^ 4);
  assign w333[20] = |(datain[231:228] ^ 0);
  assign w333[21] = |(datain[227:224] ^ 0);
  assign w333[22] = |(datain[223:220] ^ 10);
  assign w333[23] = |(datain[219:216] ^ 0);
  assign w333[24] = |(datain[215:212] ^ 1);
  assign w333[25] = |(datain[211:208] ^ 0);
  assign w333[26] = |(datain[207:204] ^ 0);
  assign w333[27] = |(datain[203:200] ^ 0);
  assign comp[333] = ~(|w333);
  wire [28-1:0] w334;
  assign w334[0] = |(datain[311:308] ^ 14);
  assign w334[1] = |(datain[307:304] ^ 15);
  assign w334[2] = |(datain[303:300] ^ 14);
  assign w334[3] = |(datain[299:296] ^ 3);
  assign w334[4] = |(datain[295:292] ^ 11);
  assign w334[5] = |(datain[291:288] ^ 15);
  assign w334[6] = |(datain[287:284] ^ 12);
  assign w334[7] = |(datain[283:280] ^ 10);
  assign w334[8] = |(datain[279:276] ^ 0);
  assign w334[9] = |(datain[275:272] ^ 3);
  assign w334[10] = |(datain[271:268] ^ 1);
  assign w334[11] = |(datain[267:264] ^ 14);
  assign w334[12] = |(datain[263:260] ^ 5);
  assign w334[13] = |(datain[259:256] ^ 7);
  assign w334[14] = |(datain[255:252] ^ 11);
  assign w334[15] = |(datain[251:248] ^ 15);
  assign w334[16] = |(datain[247:244] ^ 12);
  assign w334[17] = |(datain[243:240] ^ 10);
  assign w334[18] = |(datain[239:236] ^ 0);
  assign w334[19] = |(datain[235:232] ^ 3);
  assign w334[20] = |(datain[231:228] ^ 1);
  assign w334[21] = |(datain[227:224] ^ 14);
  assign w334[22] = |(datain[223:220] ^ 14);
  assign w334[23] = |(datain[219:216] ^ 8);
  assign w334[24] = |(datain[215:212] ^ 11);
  assign w334[25] = |(datain[211:208] ^ 4);
  assign w334[26] = |(datain[207:204] ^ 14);
  assign w334[27] = |(datain[203:200] ^ 3);
  assign comp[334] = ~(|w334);
  wire [28-1:0] w335;
  assign w335[0] = |(datain[311:308] ^ 15);
  assign w335[1] = |(datain[307:304] ^ 10);
  assign w335[2] = |(datain[303:300] ^ 11);
  assign w335[3] = |(datain[299:296] ^ 0);
  assign w335[4] = |(datain[295:292] ^ 8);
  assign w335[5] = |(datain[291:288] ^ 15);
  assign w335[6] = |(datain[287:284] ^ 5);
  assign w335[7] = |(datain[283:280] ^ 11);
  assign w335[8] = |(datain[279:276] ^ 5);
  assign w335[9] = |(datain[275:272] ^ 3);
  assign w335[10] = |(datain[271:268] ^ 11);
  assign w335[11] = |(datain[267:264] ^ 9);
  assign w335[12] = |(datain[263:260] ^ 10);
  assign w335[13] = |(datain[259:256] ^ 1);
  assign w335[14] = |(datain[255:252] ^ 0);
  assign w335[15] = |(datain[251:248] ^ 0);
  assign w335[16] = |(datain[247:244] ^ 3);
  assign w335[17] = |(datain[243:240] ^ 0);
  assign w335[18] = |(datain[239:236] ^ 0);
  assign w335[19] = |(datain[235:232] ^ 7);
  assign w335[20] = |(datain[231:228] ^ 4);
  assign w335[21] = |(datain[227:224] ^ 3);
  assign w335[22] = |(datain[223:220] ^ 14);
  assign w335[23] = |(datain[219:216] ^ 2);
  assign w335[24] = |(datain[215:212] ^ 15);
  assign w335[25] = |(datain[211:208] ^ 11);
  assign w335[26] = |(datain[207:204] ^ 12);
  assign w335[27] = |(datain[203:200] ^ 3);
  assign comp[335] = ~(|w335);
  wire [74-1:0] w336;
  assign w336[0] = |(datain[311:308] ^ 8);
  assign w336[1] = |(datain[307:304] ^ 9);
  assign w336[2] = |(datain[303:300] ^ 8);
  assign w336[3] = |(datain[299:296] ^ 6);
  assign w336[4] = |(datain[295:292] ^ 3);
  assign w336[5] = |(datain[291:288] ^ 6);
  assign w336[6] = |(datain[287:284] ^ 0);
  assign w336[7] = |(datain[283:280] ^ 1);
  assign w336[8] = |(datain[279:276] ^ 11);
  assign w336[9] = |(datain[275:272] ^ 4);
  assign w336[10] = |(datain[271:268] ^ 4);
  assign w336[11] = |(datain[267:264] ^ 0);
  assign w336[12] = |(datain[263:260] ^ 8);
  assign w336[13] = |(datain[259:256] ^ 11);
  assign w336[14] = |(datain[255:252] ^ 5);
  assign w336[15] = |(datain[251:248] ^ 14);
  assign w336[16] = |(datain[247:244] ^ 0);
  assign w336[17] = |(datain[243:240] ^ 2);
  assign w336[18] = |(datain[239:236] ^ 8);
  assign w336[19] = |(datain[235:232] ^ 13);
  assign w336[20] = |(datain[231:228] ^ 9);
  assign w336[21] = |(datain[227:224] ^ 6);
  assign w336[22] = |(datain[223:220] ^ 3);
  assign w336[23] = |(datain[219:216] ^ 5);
  assign w336[24] = |(datain[215:212] ^ 0);
  assign w336[25] = |(datain[211:208] ^ 1);
  assign w336[26] = |(datain[207:204] ^ 11);
  assign w336[27] = |(datain[203:200] ^ 9);
  assign w336[28] = |(datain[199:196] ^ 0);
  assign w336[29] = |(datain[195:192] ^ 3);
  assign w336[30] = |(datain[191:188] ^ 0);
  assign w336[31] = |(datain[187:184] ^ 0);
  assign w336[32] = |(datain[183:180] ^ 12);
  assign w336[33] = |(datain[179:176] ^ 13);
  assign w336[34] = |(datain[175:172] ^ 2);
  assign w336[35] = |(datain[171:168] ^ 1);
  assign w336[36] = |(datain[167:164] ^ 11);
  assign w336[37] = |(datain[163:160] ^ 4);
  assign w336[38] = |(datain[159:156] ^ 4);
  assign w336[39] = |(datain[155:152] ^ 2);
  assign w336[40] = |(datain[151:148] ^ 8);
  assign w336[41] = |(datain[147:144] ^ 11);
  assign w336[42] = |(datain[143:140] ^ 5);
  assign w336[43] = |(datain[139:136] ^ 14);
  assign w336[44] = |(datain[135:132] ^ 0);
  assign w336[45] = |(datain[131:128] ^ 2);
  assign w336[46] = |(datain[127:124] ^ 11);
  assign w336[47] = |(datain[123:120] ^ 9);
  assign w336[48] = |(datain[119:116] ^ 0);
  assign w336[49] = |(datain[115:112] ^ 0);
  assign w336[50] = |(datain[111:108] ^ 0);
  assign w336[51] = |(datain[107:104] ^ 0);
  assign w336[52] = |(datain[103:100] ^ 8);
  assign w336[53] = |(datain[99:96] ^ 11);
  assign w336[54] = |(datain[95:92] ^ 9);
  assign w336[55] = |(datain[91:88] ^ 6);
  assign w336[56] = |(datain[87:84] ^ 3);
  assign w336[57] = |(datain[83:80] ^ 3);
  assign w336[58] = |(datain[79:76] ^ 0);
  assign w336[59] = |(datain[75:72] ^ 1);
  assign w336[60] = |(datain[71:68] ^ 8);
  assign w336[61] = |(datain[67:64] ^ 3);
  assign w336[62] = |(datain[63:60] ^ 12);
  assign w336[63] = |(datain[59:56] ^ 2);
  assign w336[64] = |(datain[55:52] ^ 0);
  assign w336[65] = |(datain[51:48] ^ 4);
  assign w336[66] = |(datain[47:44] ^ 11);
  assign w336[67] = |(datain[43:40] ^ 0);
  assign w336[68] = |(datain[39:36] ^ 0);
  assign w336[69] = |(datain[35:32] ^ 0);
  assign w336[70] = |(datain[31:28] ^ 12);
  assign w336[71] = |(datain[27:24] ^ 13);
  assign w336[72] = |(datain[23:20] ^ 2);
  assign w336[73] = |(datain[19:16] ^ 1);
  assign comp[336] = ~(|w336);
  wire [30-1:0] w337;
  assign w337[0] = |(datain[311:308] ^ 14);
  assign w337[1] = |(datain[307:304] ^ 5);
  assign w337[2] = |(datain[303:300] ^ 8);
  assign w337[3] = |(datain[299:296] ^ 1);
  assign w337[4] = |(datain[295:292] ^ 14);
  assign w337[5] = |(datain[291:288] ^ 12);
  assign w337[6] = |(datain[287:284] ^ 0);
  assign w337[7] = |(datain[283:280] ^ 2);
  assign w337[8] = |(datain[279:276] ^ 0);
  assign w337[9] = |(datain[275:272] ^ 2);
  assign w337[10] = |(datain[271:268] ^ 11);
  assign w337[11] = |(datain[267:264] ^ 15);
  assign w337[12] = |(datain[263:260] ^ 12);
  assign w337[13] = |(datain[259:256] ^ 10);
  assign w337[14] = |(datain[255:252] ^ 0);
  assign w337[15] = |(datain[251:248] ^ 5);
  assign w337[16] = |(datain[247:244] ^ 0);
  assign w337[17] = |(datain[243:240] ^ 14);
  assign w337[18] = |(datain[239:236] ^ 5);
  assign w337[19] = |(datain[235:232] ^ 7);
  assign w337[20] = |(datain[231:228] ^ 11);
  assign w337[21] = |(datain[227:224] ^ 15);
  assign w337[22] = |(datain[223:220] ^ 3);
  assign w337[23] = |(datain[219:216] ^ 14);
  assign w337[24] = |(datain[215:212] ^ 0);
  assign w337[25] = |(datain[211:208] ^ 1);
  assign w337[26] = |(datain[207:204] ^ 1);
  assign w337[27] = |(datain[203:200] ^ 14);
  assign w337[28] = |(datain[199:196] ^ 5);
  assign w337[29] = |(datain[195:192] ^ 7);
  assign comp[337] = ~(|w337);
  wire [28-1:0] w338;
  assign w338[0] = |(datain[311:308] ^ 7);
  assign w338[1] = |(datain[307:304] ^ 5);
  assign w338[2] = |(datain[303:300] ^ 0);
  assign w338[3] = |(datain[299:296] ^ 9);
  assign w338[4] = |(datain[295:292] ^ 12);
  assign w338[5] = |(datain[291:288] ^ 4);
  assign w338[6] = |(datain[287:284] ^ 7);
  assign w338[7] = |(datain[283:280] ^ 14);
  assign w338[8] = |(datain[279:276] ^ 0);
  assign w338[9] = |(datain[275:272] ^ 4);
  assign w338[10] = |(datain[271:268] ^ 2);
  assign w338[11] = |(datain[267:264] ^ 6);
  assign w338[12] = |(datain[263:260] ^ 12);
  assign w338[13] = |(datain[259:256] ^ 6);
  assign w338[14] = |(datain[255:252] ^ 0);
  assign w338[15] = |(datain[251:248] ^ 5);
  assign w338[16] = |(datain[247:244] ^ 0);
  assign w338[17] = |(datain[243:240] ^ 0);
  assign w338[18] = |(datain[239:236] ^ 14);
  assign w338[19] = |(datain[235:232] ^ 11);
  assign w338[20] = |(datain[231:228] ^ 0);
  assign w338[21] = |(datain[227:224] ^ 15);
  assign w338[22] = |(datain[223:220] ^ 11);
  assign w338[23] = |(datain[219:216] ^ 15);
  assign w338[24] = |(datain[215:212] ^ 3);
  assign w338[25] = |(datain[211:208] ^ 15);
  assign w338[26] = |(datain[207:204] ^ 0);
  assign w338[27] = |(datain[203:200] ^ 4);
  assign comp[338] = ~(|w338);
  wire [28-1:0] w339;
  assign w339[0] = |(datain[311:308] ^ 5);
  assign w339[1] = |(datain[307:304] ^ 5);
  assign w339[2] = |(datain[303:300] ^ 8);
  assign w339[3] = |(datain[299:296] ^ 9);
  assign w339[4] = |(datain[295:292] ^ 14);
  assign w339[5] = |(datain[291:288] ^ 5);
  assign w339[6] = |(datain[287:284] ^ 8);
  assign w339[7] = |(datain[283:280] ^ 1);
  assign w339[8] = |(datain[279:276] ^ 14);
  assign w339[9] = |(datain[275:272] ^ 12);
  assign w339[10] = |(datain[271:268] ^ 0);
  assign w339[11] = |(datain[267:264] ^ 2);
  assign w339[12] = |(datain[263:260] ^ 0);
  assign w339[13] = |(datain[259:256] ^ 2);
  assign w339[14] = |(datain[255:252] ^ 11);
  assign w339[15] = |(datain[251:248] ^ 15);
  assign w339[16] = |(datain[247:244] ^ 12);
  assign w339[17] = |(datain[243:240] ^ 10);
  assign w339[18] = |(datain[239:236] ^ 0);
  assign w339[19] = |(datain[235:232] ^ 5);
  assign w339[20] = |(datain[231:228] ^ 0);
  assign w339[21] = |(datain[227:224] ^ 14);
  assign w339[22] = |(datain[223:220] ^ 5);
  assign w339[23] = |(datain[219:216] ^ 7);
  assign w339[24] = |(datain[215:212] ^ 11);
  assign w339[25] = |(datain[211:208] ^ 15);
  assign w339[26] = |(datain[207:204] ^ 3);
  assign w339[27] = |(datain[203:200] ^ 14);
  assign comp[339] = ~(|w339);
  wire [30-1:0] w340;
  assign w340[0] = |(datain[311:308] ^ 8);
  assign w340[1] = |(datain[307:304] ^ 9);
  assign w340[2] = |(datain[303:300] ^ 14);
  assign w340[3] = |(datain[299:296] ^ 5);
  assign w340[4] = |(datain[295:292] ^ 8);
  assign w340[5] = |(datain[291:288] ^ 1);
  assign w340[6] = |(datain[287:284] ^ 14);
  assign w340[7] = |(datain[283:280] ^ 12);
  assign w340[8] = |(datain[279:276] ^ 0);
  assign w340[9] = |(datain[275:272] ^ 2);
  assign w340[10] = |(datain[271:268] ^ 0);
  assign w340[11] = |(datain[267:264] ^ 2);
  assign w340[12] = |(datain[263:260] ^ 11);
  assign w340[13] = |(datain[259:256] ^ 15);
  assign w340[14] = |(datain[255:252] ^ 12);
  assign w340[15] = |(datain[251:248] ^ 10);
  assign w340[16] = |(datain[247:244] ^ 0);
  assign w340[17] = |(datain[243:240] ^ 5);
  assign w340[18] = |(datain[239:236] ^ 0);
  assign w340[19] = |(datain[235:232] ^ 14);
  assign w340[20] = |(datain[231:228] ^ 5);
  assign w340[21] = |(datain[227:224] ^ 7);
  assign w340[22] = |(datain[223:220] ^ 11);
  assign w340[23] = |(datain[219:216] ^ 15);
  assign w340[24] = |(datain[215:212] ^ 3);
  assign w340[25] = |(datain[211:208] ^ 14);
  assign w340[26] = |(datain[207:204] ^ 0);
  assign w340[27] = |(datain[203:200] ^ 1);
  assign w340[28] = |(datain[199:196] ^ 1);
  assign w340[29] = |(datain[195:192] ^ 14);
  assign comp[340] = ~(|w340);
  wire [32-1:0] w341;
  assign w341[0] = |(datain[311:308] ^ 4);
  assign w341[1] = |(datain[307:304] ^ 13);
  assign w341[2] = |(datain[303:300] ^ 5);
  assign w341[3] = |(datain[299:296] ^ 10);
  assign w341[4] = |(datain[295:292] ^ 1);
  assign w341[5] = |(datain[291:288] ^ 2);
  assign w341[6] = |(datain[287:284] ^ 0);
  assign w341[7] = |(datain[283:280] ^ 0);
  assign w341[8] = |(datain[279:276] ^ 5);
  assign w341[9] = |(datain[275:272] ^ 2);
  assign w341[10] = |(datain[271:268] ^ 0);
  assign w341[11] = |(datain[267:264] ^ 1);
  assign w341[12] = |(datain[263:260] ^ 4);
  assign w341[13] = |(datain[259:256] ^ 1);
  assign w341[14] = |(datain[255:252] ^ 1);
  assign w341[15] = |(datain[251:248] ^ 11);
  assign w341[16] = |(datain[247:244] ^ 14);
  assign w341[17] = |(datain[243:240] ^ 0);
  assign w341[18] = |(datain[239:236] ^ 0);
  assign w341[19] = |(datain[235:232] ^ 6);
  assign w341[20] = |(datain[231:228] ^ 7);
  assign w341[21] = |(datain[227:224] ^ 8);
  assign w341[22] = |(datain[223:220] ^ 0);
  assign w341[23] = |(datain[219:216] ^ 12);
  assign w341[24] = |(datain[215:212] ^ 15);
  assign w341[25] = |(datain[211:208] ^ 15);
  assign w341[26] = |(datain[207:204] ^ 15);
  assign w341[27] = |(datain[203:200] ^ 15);
  assign w341[28] = |(datain[199:196] ^ 9);
  assign w341[29] = |(datain[195:192] ^ 9);
  assign w341[30] = |(datain[191:188] ^ 2);
  assign w341[31] = |(datain[187:184] ^ 15);
  assign comp[341] = ~(|w341);
  wire [62-1:0] w342;
  assign w342[0] = |(datain[311:308] ^ 15);
  assign w342[1] = |(datain[307:304] ^ 15);
  assign w342[2] = |(datain[303:300] ^ 11);
  assign w342[3] = |(datain[299:296] ^ 14);
  assign w342[4] = |(datain[295:292] ^ 0);
  assign w342[5] = |(datain[291:288] ^ 0);
  assign w342[6] = |(datain[287:284] ^ 7);
  assign w342[7] = |(datain[283:280] ^ 12);
  assign w342[8] = |(datain[279:276] ^ 15);
  assign w342[9] = |(datain[275:272] ^ 10);
  assign w342[10] = |(datain[271:268] ^ 8);
  assign w342[11] = |(datain[267:264] ^ 11);
  assign w342[12] = |(datain[263:260] ^ 14);
  assign w342[13] = |(datain[259:256] ^ 6);
  assign w342[14] = |(datain[255:252] ^ 8);
  assign w342[15] = |(datain[251:248] ^ 14);
  assign w342[16] = |(datain[247:244] ^ 13);
  assign w342[17] = |(datain[243:240] ^ 7);
  assign w342[18] = |(datain[239:236] ^ 15);
  assign w342[19] = |(datain[235:232] ^ 11);
  assign w342[20] = |(datain[231:228] ^ 8);
  assign w342[21] = |(datain[227:224] ^ 14);
  assign w342[22] = |(datain[223:220] ^ 12);
  assign w342[23] = |(datain[219:216] ^ 7);
  assign w342[24] = |(datain[215:212] ^ 11);
  assign w342[25] = |(datain[211:208] ^ 11);
  assign w342[26] = |(datain[207:204] ^ 0);
  assign w342[27] = |(datain[203:200] ^ 0);
  assign w342[28] = |(datain[199:196] ^ 7);
  assign w342[29] = |(datain[195:192] ^ 14);
  assign w342[30] = |(datain[191:188] ^ 11);
  assign w342[31] = |(datain[187:184] ^ 8);
  assign w342[32] = |(datain[183:180] ^ 0);
  assign w342[33] = |(datain[179:176] ^ 4);
  assign w342[34] = |(datain[175:172] ^ 0);
  assign w342[35] = |(datain[171:168] ^ 2);
  assign w342[36] = |(datain[167:164] ^ 11);
  assign w342[37] = |(datain[163:160] ^ 10);
  assign w342[38] = |(datain[159:156] ^ 8);
  assign w342[39] = |(datain[155:152] ^ 0);
  assign w342[40] = |(datain[151:148] ^ 0);
  assign w342[41] = |(datain[147:144] ^ 0);
  assign w342[42] = |(datain[143:140] ^ 11);
  assign w342[43] = |(datain[139:136] ^ 9);
  assign w342[44] = |(datain[135:132] ^ 0);
  assign w342[45] = |(datain[131:128] ^ 4);
  assign w342[46] = |(datain[127:124] ^ 0);
  assign w342[47] = |(datain[123:120] ^ 0);
  assign w342[48] = |(datain[119:116] ^ 5);
  assign w342[49] = |(datain[115:112] ^ 6);
  assign w342[50] = |(datain[111:108] ^ 5);
  assign w342[51] = |(datain[107:104] ^ 3);
  assign w342[52] = |(datain[103:100] ^ 12);
  assign w342[53] = |(datain[99:96] ^ 13);
  assign w342[54] = |(datain[95:92] ^ 1);
  assign w342[55] = |(datain[91:88] ^ 3);
  assign w342[56] = |(datain[87:84] ^ 14);
  assign w342[57] = |(datain[83:80] ^ 9);
  assign w342[58] = |(datain[79:76] ^ 8);
  assign w342[59] = |(datain[75:72] ^ 0);
  assign w342[60] = |(datain[71:68] ^ 0);
  assign w342[61] = |(datain[67:64] ^ 1);
  assign comp[342] = ~(|w342);
  wire [32-1:0] w343;
  assign w343[0] = |(datain[311:308] ^ 3);
  assign w343[1] = |(datain[307:304] ^ 2);
  assign w343[2] = |(datain[303:300] ^ 14);
  assign w343[3] = |(datain[299:296] ^ 4);
  assign w343[4] = |(datain[295:292] ^ 12);
  assign w343[5] = |(datain[291:288] ^ 13);
  assign w343[6] = |(datain[287:284] ^ 1);
  assign w343[7] = |(datain[283:280] ^ 6);
  assign w343[8] = |(datain[279:276] ^ 12);
  assign w343[9] = |(datain[275:272] ^ 13);
  assign w343[10] = |(datain[271:268] ^ 1);
  assign w343[11] = |(datain[267:264] ^ 2);
  assign w343[12] = |(datain[263:260] ^ 3);
  assign w343[13] = |(datain[259:256] ^ 3);
  assign w343[14] = |(datain[255:252] ^ 12);
  assign w343[15] = |(datain[251:248] ^ 0);
  assign w343[16] = |(datain[247:244] ^ 12);
  assign w343[17] = |(datain[243:240] ^ 13);
  assign w343[18] = |(datain[239:236] ^ 1);
  assign w343[19] = |(datain[235:232] ^ 3);
  assign w343[20] = |(datain[231:228] ^ 0);
  assign w343[21] = |(datain[227:224] ^ 14);
  assign w343[22] = |(datain[223:220] ^ 0);
  assign w343[23] = |(datain[219:216] ^ 7);
  assign w343[24] = |(datain[215:212] ^ 11);
  assign w343[25] = |(datain[211:208] ^ 8);
  assign w343[26] = |(datain[207:204] ^ 0);
  assign w343[27] = |(datain[203:200] ^ 0);
  assign w343[28] = |(datain[199:196] ^ 0);
  assign w343[29] = |(datain[195:192] ^ 2);
  assign w343[30] = |(datain[191:188] ^ 11);
  assign w343[31] = |(datain[187:184] ^ 9);
  assign comp[343] = ~(|w343);
  wire [30-1:0] w344;
  assign w344[0] = |(datain[311:308] ^ 10);
  assign w344[1] = |(datain[307:304] ^ 3);
  assign w344[2] = |(datain[303:300] ^ 11);
  assign w344[3] = |(datain[299:296] ^ 8);
  assign w344[4] = |(datain[295:292] ^ 7);
  assign w344[5] = |(datain[291:288] ^ 13);
  assign w344[6] = |(datain[287:284] ^ 11);
  assign w344[7] = |(datain[283:280] ^ 8);
  assign w344[8] = |(datain[279:276] ^ 3);
  assign w344[9] = |(datain[275:272] ^ 1);
  assign w344[10] = |(datain[271:268] ^ 0);
  assign w344[11] = |(datain[267:264] ^ 1);
  assign w344[12] = |(datain[263:260] ^ 10);
  assign w344[13] = |(datain[259:256] ^ 3);
  assign w344[14] = |(datain[255:252] ^ 11);
  assign w344[15] = |(datain[251:248] ^ 12);
  assign w344[16] = |(datain[247:244] ^ 7);
  assign w344[17] = |(datain[243:240] ^ 13);
  assign w344[18] = |(datain[239:236] ^ 15);
  assign w344[19] = |(datain[235:232] ^ 15);
  assign w344[20] = |(datain[231:228] ^ 0);
  assign w344[21] = |(datain[227:224] ^ 14);
  assign w344[22] = |(datain[223:220] ^ 1);
  assign w344[23] = |(datain[219:216] ^ 3);
  assign w344[24] = |(datain[215:212] ^ 0);
  assign w344[25] = |(datain[211:208] ^ 4);
  assign w344[26] = |(datain[207:204] ^ 12);
  assign w344[27] = |(datain[203:200] ^ 13);
  assign w344[28] = |(datain[199:196] ^ 1);
  assign w344[29] = |(datain[195:192] ^ 2);
  assign comp[344] = ~(|w344);
  wire [38-1:0] w345;
  assign w345[0] = |(datain[311:308] ^ 1);
  assign w345[1] = |(datain[307:304] ^ 14);
  assign w345[2] = |(datain[303:300] ^ 5);
  assign w345[3] = |(datain[299:296] ^ 3);
  assign w345[4] = |(datain[295:292] ^ 15);
  assign w345[5] = |(datain[291:288] ^ 15);
  assign w345[6] = |(datain[287:284] ^ 0);
  assign w345[7] = |(datain[283:280] ^ 14);
  assign w345[8] = |(datain[279:276] ^ 1);
  assign w345[9] = |(datain[275:272] ^ 3);
  assign w345[10] = |(datain[271:268] ^ 0);
  assign w345[11] = |(datain[267:264] ^ 4);
  assign w345[12] = |(datain[263:260] ^ 12);
  assign w345[13] = |(datain[259:256] ^ 13);
  assign w345[14] = |(datain[255:252] ^ 1);
  assign w345[15] = |(datain[251:248] ^ 2);
  assign w345[16] = |(datain[247:244] ^ 11);
  assign w345[17] = |(datain[243:240] ^ 1);
  assign w345[18] = |(datain[239:236] ^ 0);
  assign w345[19] = |(datain[235:232] ^ 6);
  assign w345[20] = |(datain[231:228] ^ 13);
  assign w345[21] = |(datain[227:224] ^ 3);
  assign w345[22] = |(datain[223:220] ^ 14);
  assign w345[23] = |(datain[219:216] ^ 0);
  assign w345[24] = |(datain[215:212] ^ 8);
  assign w345[25] = |(datain[211:208] ^ 14);
  assign w345[26] = |(datain[207:204] ^ 12);
  assign w345[27] = |(datain[203:200] ^ 0);
  assign w345[28] = |(datain[199:196] ^ 8);
  assign w345[29] = |(datain[195:192] ^ 7);
  assign w345[30] = |(datain[191:188] ^ 0);
  assign w345[31] = |(datain[187:184] ^ 6);
  assign w345[32] = |(datain[183:180] ^ 4);
  assign w345[33] = |(datain[179:176] ^ 14);
  assign w345[34] = |(datain[175:172] ^ 0);
  assign w345[35] = |(datain[171:168] ^ 0);
  assign w345[36] = |(datain[167:164] ^ 10);
  assign w345[37] = |(datain[163:160] ^ 3);
  assign comp[345] = ~(|w345);
  wire [28-1:0] w346;
  assign w346[0] = |(datain[311:308] ^ 12);
  assign w346[1] = |(datain[307:304] ^ 13);
  assign w346[2] = |(datain[303:300] ^ 1);
  assign w346[3] = |(datain[299:296] ^ 6);
  assign w346[4] = |(datain[295:292] ^ 3);
  assign w346[5] = |(datain[291:288] ^ 3);
  assign w346[6] = |(datain[287:284] ^ 12);
  assign w346[7] = |(datain[283:280] ^ 0);
  assign w346[8] = |(datain[279:276] ^ 12);
  assign w346[9] = |(datain[275:272] ^ 13);
  assign w346[10] = |(datain[271:268] ^ 1);
  assign w346[11] = |(datain[267:264] ^ 3);
  assign w346[12] = |(datain[263:260] ^ 0);
  assign w346[13] = |(datain[259:256] ^ 14);
  assign w346[14] = |(datain[255:252] ^ 0);
  assign w346[15] = |(datain[251:248] ^ 7);
  assign w346[16] = |(datain[247:244] ^ 11);
  assign w346[17] = |(datain[243:240] ^ 11);
  assign w346[18] = |(datain[239:236] ^ 0);
  assign w346[19] = |(datain[235:232] ^ 0);
  assign w346[20] = |(datain[231:228] ^ 0);
  assign w346[21] = |(datain[227:224] ^ 2);
  assign w346[22] = |(datain[223:220] ^ 11);
  assign w346[23] = |(datain[219:216] ^ 9);
  assign w346[24] = |(datain[215:212] ^ 0);
  assign w346[25] = |(datain[211:208] ^ 6);
  assign w346[26] = |(datain[207:204] ^ 0);
  assign w346[27] = |(datain[203:200] ^ 0);
  assign comp[346] = ~(|w346);
  wire [32-1:0] w347;
  assign w347[0] = |(datain[311:308] ^ 3);
  assign w347[1] = |(datain[307:304] ^ 2);
  assign w347[2] = |(datain[303:300] ^ 14);
  assign w347[3] = |(datain[299:296] ^ 4);
  assign w347[4] = |(datain[295:292] ^ 12);
  assign w347[5] = |(datain[291:288] ^ 13);
  assign w347[6] = |(datain[287:284] ^ 1);
  assign w347[7] = |(datain[283:280] ^ 6);
  assign w347[8] = |(datain[279:276] ^ 12);
  assign w347[9] = |(datain[275:272] ^ 13);
  assign w347[10] = |(datain[271:268] ^ 1);
  assign w347[11] = |(datain[267:264] ^ 2);
  assign w347[12] = |(datain[263:260] ^ 3);
  assign w347[13] = |(datain[259:256] ^ 3);
  assign w347[14] = |(datain[255:252] ^ 12);
  assign w347[15] = |(datain[251:248] ^ 0);
  assign w347[16] = |(datain[247:244] ^ 12);
  assign w347[17] = |(datain[243:240] ^ 13);
  assign w347[18] = |(datain[239:236] ^ 1);
  assign w347[19] = |(datain[235:232] ^ 3);
  assign w347[20] = |(datain[231:228] ^ 0);
  assign w347[21] = |(datain[227:224] ^ 14);
  assign w347[22] = |(datain[223:220] ^ 0);
  assign w347[23] = |(datain[219:216] ^ 7);
  assign w347[24] = |(datain[215:212] ^ 11);
  assign w347[25] = |(datain[211:208] ^ 11);
  assign w347[26] = |(datain[207:204] ^ 0);
  assign w347[27] = |(datain[203:200] ^ 0);
  assign w347[28] = |(datain[199:196] ^ 0);
  assign w347[29] = |(datain[195:192] ^ 2);
  assign w347[30] = |(datain[191:188] ^ 11);
  assign w347[31] = |(datain[187:184] ^ 9);
  assign comp[347] = ~(|w347);
  wire [30-1:0] w348;
  assign w348[0] = |(datain[311:308] ^ 12);
  assign w348[1] = |(datain[307:304] ^ 4);
  assign w348[2] = |(datain[303:300] ^ 7);
  assign w348[3] = |(datain[299:296] ^ 13);
  assign w348[4] = |(datain[295:292] ^ 11);
  assign w348[5] = |(datain[291:288] ^ 8);
  assign w348[6] = |(datain[287:284] ^ 14);
  assign w348[7] = |(datain[283:280] ^ 4);
  assign w348[8] = |(datain[279:276] ^ 0);
  assign w348[9] = |(datain[275:272] ^ 0);
  assign w348[10] = |(datain[271:268] ^ 10);
  assign w348[11] = |(datain[267:264] ^ 3);
  assign w348[12] = |(datain[263:260] ^ 11);
  assign w348[13] = |(datain[259:256] ^ 8);
  assign w348[14] = |(datain[255:252] ^ 7);
  assign w348[15] = |(datain[251:248] ^ 13);
  assign w348[16] = |(datain[247:244] ^ 11);
  assign w348[17] = |(datain[243:240] ^ 8);
  assign w348[18] = |(datain[239:236] ^ 3);
  assign w348[19] = |(datain[235:232] ^ 1);
  assign w348[20] = |(datain[231:228] ^ 0);
  assign w348[21] = |(datain[227:224] ^ 1);
  assign w348[22] = |(datain[223:220] ^ 10);
  assign w348[23] = |(datain[219:216] ^ 3);
  assign w348[24] = |(datain[215:212] ^ 11);
  assign w348[25] = |(datain[211:208] ^ 12);
  assign w348[26] = |(datain[207:204] ^ 7);
  assign w348[27] = |(datain[203:200] ^ 13);
  assign w348[28] = |(datain[199:196] ^ 15);
  assign w348[29] = |(datain[195:192] ^ 15);
  assign comp[348] = ~(|w348);
  wire [36-1:0] w349;
  assign w349[0] = |(datain[311:308] ^ 2);
  assign w349[1] = |(datain[307:304] ^ 14);
  assign w349[2] = |(datain[303:300] ^ 12);
  assign w349[3] = |(datain[299:296] ^ 0);
  assign w349[4] = |(datain[295:292] ^ 0);
  assign w349[5] = |(datain[291:288] ^ 1);
  assign w349[6] = |(datain[287:284] ^ 5);
  assign w349[7] = |(datain[283:280] ^ 3);
  assign w349[8] = |(datain[279:276] ^ 0);
  assign w349[9] = |(datain[275:272] ^ 14);
  assign w349[10] = |(datain[271:268] ^ 14);
  assign w349[11] = |(datain[267:264] ^ 8);
  assign w349[12] = |(datain[263:260] ^ 11);
  assign w349[13] = |(datain[259:256] ^ 1);
  assign w349[14] = |(datain[255:252] ^ 15);
  assign w349[15] = |(datain[251:248] ^ 15);
  assign w349[16] = |(datain[247:244] ^ 0);
  assign w349[17] = |(datain[243:240] ^ 14);
  assign w349[18] = |(datain[239:236] ^ 11);
  assign w349[19] = |(datain[235:232] ^ 11);
  assign w349[20] = |(datain[231:228] ^ 4);
  assign w349[21] = |(datain[227:224] ^ 12);
  assign w349[22] = |(datain[223:220] ^ 0);
  assign w349[23] = |(datain[219:216] ^ 0);
  assign w349[24] = |(datain[215:212] ^ 14);
  assign w349[25] = |(datain[211:208] ^ 8);
  assign w349[26] = |(datain[207:204] ^ 10);
  assign w349[27] = |(datain[203:200] ^ 13);
  assign w349[28] = |(datain[199:196] ^ 15);
  assign w349[29] = |(datain[195:192] ^ 15);
  assign w349[30] = |(datain[191:188] ^ 5);
  assign w349[31] = |(datain[187:184] ^ 11);
  assign w349[32] = |(datain[183:180] ^ 12);
  assign w349[33] = |(datain[179:176] ^ 13);
  assign w349[34] = |(datain[175:172] ^ 1);
  assign w349[35] = |(datain[171:168] ^ 2);
  assign comp[349] = ~(|w349);
  wire [46-1:0] w350;
  assign w350[0] = |(datain[311:308] ^ 7);
  assign w350[1] = |(datain[307:304] ^ 2);
  assign w350[2] = |(datain[303:300] ^ 6);
  assign w350[3] = |(datain[299:296] ^ 1);
  assign w350[4] = |(datain[295:292] ^ 12);
  assign w350[5] = |(datain[291:288] ^ 13);
  assign w350[6] = |(datain[287:284] ^ 2);
  assign w350[7] = |(datain[283:280] ^ 1);
  assign w350[8] = |(datain[279:276] ^ 0);
  assign w350[9] = |(datain[275:272] ^ 10);
  assign w350[10] = |(datain[271:268] ^ 12);
  assign w350[11] = |(datain[267:264] ^ 0);
  assign w350[12] = |(datain[263:260] ^ 7);
  assign w350[13] = |(datain[259:256] ^ 5);
  assign w350[14] = |(datain[255:252] ^ 4);
  assign w350[15] = |(datain[251:248] ^ 12);
  assign w350[16] = |(datain[247:244] ^ 5);
  assign w350[17] = |(datain[243:240] ^ 6);
  assign w350[18] = |(datain[239:236] ^ 3);
  assign w350[19] = |(datain[235:232] ^ 3);
  assign w350[20] = |(datain[231:228] ^ 15);
  assign w350[21] = |(datain[227:224] ^ 15);
  assign w350[22] = |(datain[223:220] ^ 1);
  assign w350[23] = |(datain[219:216] ^ 14);
  assign w350[24] = |(datain[215:212] ^ 8);
  assign w350[25] = |(datain[211:208] ^ 12);
  assign w350[26] = |(datain[207:204] ^ 12);
  assign w350[27] = |(datain[203:200] ^ 8);
  assign w350[28] = |(datain[199:196] ^ 4);
  assign w350[29] = |(datain[195:192] ^ 8);
  assign w350[30] = |(datain[191:188] ^ 8);
  assign w350[31] = |(datain[187:184] ^ 14);
  assign w350[32] = |(datain[183:180] ^ 13);
  assign w350[33] = |(datain[179:176] ^ 8);
  assign w350[34] = |(datain[175:172] ^ 11);
  assign w350[35] = |(datain[171:168] ^ 11);
  assign w350[36] = |(datain[167:164] ^ 1);
  assign w350[37] = |(datain[163:160] ^ 10);
  assign w350[38] = |(datain[159:156] ^ 0);
  assign w350[39] = |(datain[155:152] ^ 0);
  assign w350[40] = |(datain[151:148] ^ 12);
  assign w350[41] = |(datain[147:144] ^ 6);
  assign w350[42] = |(datain[143:140] ^ 0);
  assign w350[43] = |(datain[139:136] ^ 5);
  assign w350[44] = |(datain[135:132] ^ 4);
  assign w350[45] = |(datain[131:128] ^ 13);
  assign comp[350] = ~(|w350);
  wire [46-1:0] w351;
  assign w351[0] = |(datain[311:308] ^ 6);
  assign w351[1] = |(datain[307:304] ^ 7);
  assign w351[2] = |(datain[303:300] ^ 0);
  assign w351[3] = |(datain[299:296] ^ 0);
  assign w351[4] = |(datain[295:292] ^ 15);
  assign w351[5] = |(datain[291:288] ^ 8);
  assign w351[6] = |(datain[287:284] ^ 11);
  assign w351[7] = |(datain[283:280] ^ 8);
  assign w351[8] = |(datain[279:276] ^ 10);
  assign w351[9] = |(datain[275:272] ^ 13);
  assign w351[10] = |(datain[271:268] ^ 13);
  assign w351[11] = |(datain[267:264] ^ 14);
  assign w351[12] = |(datain[263:260] ^ 12);
  assign w351[13] = |(datain[259:256] ^ 13);
  assign w351[14] = |(datain[255:252] ^ 2);
  assign w351[15] = |(datain[251:248] ^ 1);
  assign w351[16] = |(datain[247:244] ^ 7);
  assign w351[17] = |(datain[243:240] ^ 2);
  assign w351[18] = |(datain[239:236] ^ 4);
  assign w351[19] = |(datain[235:232] ^ 11);
  assign w351[20] = |(datain[231:228] ^ 14);
  assign w351[21] = |(datain[227:224] ^ 8);
  assign w351[22] = |(datain[223:220] ^ 7);
  assign w351[23] = |(datain[219:216] ^ 4);
  assign w351[24] = |(datain[215:212] ^ 0);
  assign w351[25] = |(datain[211:208] ^ 2);
  assign w351[26] = |(datain[207:204] ^ 0);
  assign w351[27] = |(datain[203:200] ^ 14);
  assign w351[28] = |(datain[199:196] ^ 0);
  assign w351[29] = |(datain[195:192] ^ 7);
  assign w351[30] = |(datain[191:188] ^ 3);
  assign w351[31] = |(datain[187:184] ^ 2);
  assign w351[32] = |(datain[183:180] ^ 12);
  assign w351[33] = |(datain[179:176] ^ 0);
  assign w351[34] = |(datain[175:172] ^ 11);
  assign w351[35] = |(datain[171:168] ^ 9);
  assign w351[36] = |(datain[167:164] ^ 1);
  assign w351[37] = |(datain[163:160] ^ 12);
  assign w351[38] = |(datain[159:156] ^ 0);
  assign w351[39] = |(datain[155:152] ^ 0);
  assign w351[40] = |(datain[151:148] ^ 11);
  assign w351[41] = |(datain[147:144] ^ 15);
  assign w351[42] = |(datain[143:140] ^ 10);
  assign w351[43] = |(datain[139:136] ^ 6);
  assign w351[44] = |(datain[135:132] ^ 0);
  assign w351[45] = |(datain[131:128] ^ 2);
  assign comp[351] = ~(|w351);
  wire [42-1:0] w352;
  assign w352[0] = |(datain[311:308] ^ 12);
  assign w352[1] = |(datain[307:304] ^ 13);
  assign w352[2] = |(datain[303:300] ^ 2);
  assign w352[3] = |(datain[299:296] ^ 1);
  assign w352[4] = |(datain[295:292] ^ 7);
  assign w352[5] = |(datain[291:288] ^ 2);
  assign w352[6] = |(datain[287:284] ^ 4);
  assign w352[7] = |(datain[283:280] ^ 11);
  assign w352[8] = |(datain[279:276] ^ 14);
  assign w352[9] = |(datain[275:272] ^ 8);
  assign w352[10] = |(datain[271:268] ^ 2);
  assign w352[11] = |(datain[267:264] ^ 2);
  assign w352[12] = |(datain[263:260] ^ 0);
  assign w352[13] = |(datain[259:256] ^ 3);
  assign w352[14] = |(datain[255:252] ^ 0);
  assign w352[15] = |(datain[251:248] ^ 14);
  assign w352[16] = |(datain[247:244] ^ 0);
  assign w352[17] = |(datain[243:240] ^ 7);
  assign w352[18] = |(datain[239:236] ^ 3);
  assign w352[19] = |(datain[235:232] ^ 2);
  assign w352[20] = |(datain[231:228] ^ 12);
  assign w352[21] = |(datain[227:224] ^ 0);
  assign w352[22] = |(datain[223:220] ^ 11);
  assign w352[23] = |(datain[219:216] ^ 9);
  assign w352[24] = |(datain[215:212] ^ 6);
  assign w352[25] = |(datain[211:208] ^ 13);
  assign w352[26] = |(datain[207:204] ^ 0);
  assign w352[27] = |(datain[203:200] ^ 0);
  assign w352[28] = |(datain[199:196] ^ 11);
  assign w352[29] = |(datain[195:192] ^ 15);
  assign w352[30] = |(datain[191:188] ^ 5);
  assign w352[31] = |(datain[187:184] ^ 4);
  assign w352[32] = |(datain[183:180] ^ 0);
  assign w352[33] = |(datain[179:176] ^ 3);
  assign w352[34] = |(datain[175:172] ^ 15);
  assign w352[35] = |(datain[171:168] ^ 12);
  assign w352[36] = |(datain[167:164] ^ 15);
  assign w352[37] = |(datain[163:160] ^ 3);
  assign w352[38] = |(datain[159:156] ^ 10);
  assign w352[39] = |(datain[155:152] ^ 10);
  assign w352[40] = |(datain[151:148] ^ 8);
  assign w352[41] = |(datain[147:144] ^ 12);
  assign comp[352] = ~(|w352);
  wire [74-1:0] w353;
  assign w353[0] = |(datain[311:308] ^ 0);
  assign w353[1] = |(datain[307:304] ^ 1);
  assign w353[2] = |(datain[303:300] ^ 4);
  assign w353[3] = |(datain[299:296] ^ 1);
  assign w353[4] = |(datain[295:292] ^ 4);
  assign w353[5] = |(datain[291:288] ^ 10);
  assign w353[6] = |(datain[287:284] ^ 8);
  assign w353[7] = |(datain[283:280] ^ 3);
  assign w353[8] = |(datain[279:276] ^ 0);
  assign w353[9] = |(datain[275:272] ^ 6);
  assign w353[10] = |(datain[271:268] ^ 7);
  assign w353[11] = |(datain[267:264] ^ 0);
  assign w353[12] = |(datain[263:260] ^ 0);
  assign w353[13] = |(datain[259:256] ^ 1);
  assign w353[14] = |(datain[255:252] ^ 2);
  assign w353[15] = |(datain[251:248] ^ 9);
  assign w353[16] = |(datain[247:244] ^ 11);
  assign w353[17] = |(datain[243:240] ^ 8);
  assign w353[18] = |(datain[239:236] ^ 0);
  assign w353[19] = |(datain[235:232] ^ 0);
  assign w353[20] = |(datain[231:228] ^ 4);
  assign w353[21] = |(datain[227:224] ^ 2);
  assign w353[22] = |(datain[223:220] ^ 9);
  assign w353[23] = |(datain[219:216] ^ 9);
  assign w353[24] = |(datain[215:212] ^ 3);
  assign w353[25] = |(datain[211:208] ^ 3);
  assign w353[26] = |(datain[207:204] ^ 12);
  assign w353[27] = |(datain[203:200] ^ 9);
  assign w353[28] = |(datain[199:196] ^ 12);
  assign w353[29] = |(datain[195:192] ^ 13);
  assign w353[30] = |(datain[191:188] ^ 2);
  assign w353[31] = |(datain[187:184] ^ 1);
  assign w353[32] = |(datain[183:180] ^ 11);
  assign w353[33] = |(datain[179:176] ^ 4);
  assign w353[34] = |(datain[175:172] ^ 4);
  assign w353[35] = |(datain[171:168] ^ 0);
  assign w353[36] = |(datain[167:164] ^ 11);
  assign w353[37] = |(datain[163:160] ^ 9);
  assign w353[38] = |(datain[159:156] ^ 2);
  assign w353[39] = |(datain[155:152] ^ 0);
  assign w353[40] = |(datain[151:148] ^ 0);
  assign w353[41] = |(datain[147:144] ^ 0);
  assign w353[42] = |(datain[143:140] ^ 11);
  assign w353[43] = |(datain[139:136] ^ 10);
  assign w353[44] = |(datain[135:132] ^ 6);
  assign w353[45] = |(datain[131:128] ^ 6);
  assign w353[46] = |(datain[127:124] ^ 0);
  assign w353[47] = |(datain[123:120] ^ 1);
  assign w353[48] = |(datain[119:116] ^ 12);
  assign w353[49] = |(datain[115:112] ^ 13);
  assign w353[50] = |(datain[111:108] ^ 2);
  assign w353[51] = |(datain[107:104] ^ 1);
  assign w353[52] = |(datain[103:100] ^ 11);
  assign w353[53] = |(datain[99:96] ^ 4);
  assign w353[54] = |(datain[95:92] ^ 0);
  assign w353[55] = |(datain[91:88] ^ 2);
  assign w353[56] = |(datain[87:84] ^ 11);
  assign w353[57] = |(datain[83:80] ^ 2);
  assign w353[58] = |(datain[79:76] ^ 0);
  assign w353[59] = |(datain[75:72] ^ 7);
  assign w353[60] = |(datain[71:68] ^ 12);
  assign w353[61] = |(datain[67:64] ^ 13);
  assign w353[62] = |(datain[63:60] ^ 2);
  assign w353[63] = |(datain[59:56] ^ 1);
  assign w353[64] = |(datain[55:52] ^ 11);
  assign w353[65] = |(datain[51:48] ^ 4);
  assign w353[66] = |(datain[47:44] ^ 3);
  assign w353[67] = |(datain[43:40] ^ 14);
  assign w353[68] = |(datain[39:36] ^ 12);
  assign w353[69] = |(datain[35:32] ^ 13);
  assign w353[70] = |(datain[31:28] ^ 2);
  assign w353[71] = |(datain[27:24] ^ 1);
  assign w353[72] = |(datain[23:20] ^ 1);
  assign w353[73] = |(datain[19:16] ^ 15);
  assign comp[353] = ~(|w353);
  wire [74-1:0] w354;
  assign w354[0] = |(datain[311:308] ^ 7);
  assign w354[1] = |(datain[307:304] ^ 7);
  assign w354[2] = |(datain[303:300] ^ 11);
  assign w354[3] = |(datain[299:296] ^ 1);
  assign w354[4] = |(datain[295:292] ^ 3);
  assign w354[5] = |(datain[291:288] ^ 14);
  assign w354[6] = |(datain[287:284] ^ 8);
  assign w354[7] = |(datain[283:280] ^ 9);
  assign w354[8] = |(datain[279:276] ^ 8);
  assign w354[9] = |(datain[275:272] ^ 6);
  assign w354[10] = |(datain[271:268] ^ 15);
  assign w354[11] = |(datain[267:264] ^ 14);
  assign w354[12] = |(datain[263:260] ^ 0);
  assign w354[13] = |(datain[259:256] ^ 1);
  assign w354[14] = |(datain[255:252] ^ 2);
  assign w354[15] = |(datain[251:248] ^ 13);
  assign w354[16] = |(datain[247:244] ^ 0);
  assign w354[17] = |(datain[243:240] ^ 3);
  assign w354[18] = |(datain[239:236] ^ 0);
  assign w354[19] = |(datain[235:232] ^ 0);
  assign w354[20] = |(datain[231:228] ^ 2);
  assign w354[21] = |(datain[227:224] ^ 14);
  assign w354[22] = |(datain[223:220] ^ 8);
  assign w354[23] = |(datain[219:216] ^ 9);
  assign w354[24] = |(datain[215:212] ^ 8);
  assign w354[25] = |(datain[211:208] ^ 6);
  assign w354[26] = |(datain[207:204] ^ 15);
  assign w354[27] = |(datain[203:200] ^ 3);
  assign w354[28] = |(datain[199:196] ^ 0);
  assign w354[29] = |(datain[195:192] ^ 0);
  assign w354[30] = |(datain[191:188] ^ 11);
  assign w354[31] = |(datain[187:184] ^ 8);
  assign w354[32] = |(datain[183:180] ^ 0);
  assign w354[33] = |(datain[179:176] ^ 0);
  assign w354[34] = |(datain[175:172] ^ 4);
  assign w354[35] = |(datain[171:168] ^ 2);
  assign w354[36] = |(datain[167:164] ^ 3);
  assign w354[37] = |(datain[163:160] ^ 3);
  assign w354[38] = |(datain[159:156] ^ 12);
  assign w354[39] = |(datain[155:152] ^ 9);
  assign w354[40] = |(datain[151:148] ^ 3);
  assign w354[41] = |(datain[147:144] ^ 3);
  assign w354[42] = |(datain[143:140] ^ 13);
  assign w354[43] = |(datain[139:136] ^ 2);
  assign w354[44] = |(datain[135:132] ^ 12);
  assign w354[45] = |(datain[131:128] ^ 13);
  assign w354[46] = |(datain[127:124] ^ 2);
  assign w354[47] = |(datain[123:120] ^ 1);
  assign w354[48] = |(datain[119:116] ^ 11);
  assign w354[49] = |(datain[115:112] ^ 4);
  assign w354[50] = |(datain[111:108] ^ 4);
  assign w354[51] = |(datain[107:104] ^ 0);
  assign w354[52] = |(datain[103:100] ^ 11);
  assign w354[53] = |(datain[99:96] ^ 9);
  assign w354[54] = |(datain[95:92] ^ 0);
  assign w354[55] = |(datain[91:88] ^ 5);
  assign w354[56] = |(datain[87:84] ^ 0);
  assign w354[57] = |(datain[83:80] ^ 0);
  assign w354[58] = |(datain[79:76] ^ 8);
  assign w354[59] = |(datain[75:72] ^ 11);
  assign w354[60] = |(datain[71:68] ^ 13);
  assign w354[61] = |(datain[67:64] ^ 5);
  assign w354[62] = |(datain[63:60] ^ 8);
  assign w354[63] = |(datain[59:56] ^ 1);
  assign w354[64] = |(datain[55:52] ^ 12);
  assign w354[65] = |(datain[51:48] ^ 2);
  assign w354[66] = |(datain[47:44] ^ 15);
  assign w354[67] = |(datain[43:40] ^ 2);
  assign w354[68] = |(datain[39:36] ^ 0);
  assign w354[69] = |(datain[35:32] ^ 0);
  assign w354[70] = |(datain[31:28] ^ 12);
  assign w354[71] = |(datain[27:24] ^ 13);
  assign w354[72] = |(datain[23:20] ^ 2);
  assign w354[73] = |(datain[19:16] ^ 1);
  assign comp[354] = ~(|w354);
  wire [32-1:0] w355;
  assign w355[0] = |(datain[311:308] ^ 14);
  assign w355[1] = |(datain[307:304] ^ 8);
  assign w355[2] = |(datain[303:300] ^ 0);
  assign w355[3] = |(datain[299:296] ^ 0);
  assign w355[4] = |(datain[295:292] ^ 0);
  assign w355[5] = |(datain[291:288] ^ 0);
  assign w355[6] = |(datain[287:284] ^ 5);
  assign w355[7] = |(datain[283:280] ^ 14);
  assign w355[8] = |(datain[279:276] ^ 8);
  assign w355[9] = |(datain[275:272] ^ 11);
  assign w355[10] = |(datain[271:268] ^ 13);
  assign w355[11] = |(datain[267:264] ^ 6);
  assign w355[12] = |(datain[263:260] ^ 8);
  assign w355[13] = |(datain[259:256] ^ 1);
  assign w355[14] = |(datain[255:252] ^ 12);
  assign w355[15] = |(datain[251:248] ^ 6);
  assign w355[16] = |(datain[247:244] ^ 2);
  assign w355[17] = |(datain[243:240] ^ 10);
  assign w355[18] = |(datain[239:236] ^ 0);
  assign w355[19] = |(datain[235:232] ^ 1);
  assign w355[20] = |(datain[231:228] ^ 11);
  assign w355[21] = |(datain[227:224] ^ 15);
  assign w355[22] = |(datain[223:220] ^ 0);
  assign w355[23] = |(datain[219:216] ^ 0);
  assign w355[24] = |(datain[215:212] ^ 0);
  assign w355[25] = |(datain[211:208] ^ 1);
  assign w355[26] = |(datain[207:204] ^ 10);
  assign w355[27] = |(datain[203:200] ^ 5);
  assign w355[28] = |(datain[199:196] ^ 10);
  assign w355[29] = |(datain[195:192] ^ 4);
  assign w355[30] = |(datain[191:188] ^ 8);
  assign w355[31] = |(datain[187:184] ^ 1);
  assign comp[355] = ~(|w355);
  wire [34-1:0] w356;
  assign w356[0] = |(datain[311:308] ^ 4);
  assign w356[1] = |(datain[307:304] ^ 0);
  assign w356[2] = |(datain[303:300] ^ 12);
  assign w356[3] = |(datain[299:296] ^ 13);
  assign w356[4] = |(datain[295:292] ^ 2);
  assign w356[5] = |(datain[291:288] ^ 1);
  assign w356[6] = |(datain[287:284] ^ 7);
  assign w356[7] = |(datain[283:280] ^ 2);
  assign w356[8] = |(datain[279:276] ^ 6);
  assign w356[9] = |(datain[275:272] ^ 0);
  assign w356[10] = |(datain[271:268] ^ 8);
  assign w356[11] = |(datain[267:264] ^ 11);
  assign w356[12] = |(datain[263:260] ^ 13);
  assign w356[13] = |(datain[259:256] ^ 6);
  assign w356[14] = |(datain[255:252] ^ 8);
  assign w356[15] = |(datain[251:248] ^ 3);
  assign w356[16] = |(datain[247:244] ^ 12);
  assign w356[17] = |(datain[243:240] ^ 2);
  assign w356[18] = |(datain[239:236] ^ 1);
  assign w356[19] = |(datain[235:232] ^ 4);
  assign w356[20] = |(datain[231:228] ^ 11);
  assign w356[21] = |(datain[227:224] ^ 4);
  assign w356[22] = |(datain[223:220] ^ 4);
  assign w356[23] = |(datain[219:216] ^ 0);
  assign w356[24] = |(datain[215:212] ^ 11);
  assign w356[25] = |(datain[211:208] ^ 9);
  assign w356[26] = |(datain[207:204] ^ 0);
  assign w356[27] = |(datain[203:200] ^ 4);
  assign w356[28] = |(datain[199:196] ^ 0);
  assign w356[29] = |(datain[195:192] ^ 0);
  assign w356[30] = |(datain[191:188] ^ 12);
  assign w356[31] = |(datain[187:184] ^ 13);
  assign w356[32] = |(datain[183:180] ^ 2);
  assign w356[33] = |(datain[179:176] ^ 1);
  assign comp[356] = ~(|w356);
  wire [44-1:0] w357;
  assign w357[0] = |(datain[311:308] ^ 0);
  assign w357[1] = |(datain[307:304] ^ 1);
  assign w357[2] = |(datain[303:300] ^ 0);
  assign w357[3] = |(datain[299:296] ^ 3);
  assign w357[4] = |(datain[295:292] ^ 13);
  assign w357[5] = |(datain[291:288] ^ 6);
  assign w357[6] = |(datain[287:284] ^ 11);
  assign w357[7] = |(datain[283:280] ^ 4);
  assign w357[8] = |(datain[279:276] ^ 4);
  assign w357[9] = |(datain[275:272] ^ 0);
  assign w357[10] = |(datain[271:268] ^ 12);
  assign w357[11] = |(datain[267:264] ^ 13);
  assign w357[12] = |(datain[263:260] ^ 2);
  assign w357[13] = |(datain[259:256] ^ 1);
  assign w357[14] = |(datain[255:252] ^ 3);
  assign w357[15] = |(datain[251:248] ^ 3);
  assign w357[16] = |(datain[247:244] ^ 12);
  assign w357[17] = |(datain[243:240] ^ 9);
  assign w357[18] = |(datain[239:236] ^ 3);
  assign w357[19] = |(datain[235:232] ^ 3);
  assign w357[20] = |(datain[231:228] ^ 13);
  assign w357[21] = |(datain[227:224] ^ 2);
  assign w357[22] = |(datain[223:220] ^ 3);
  assign w357[23] = |(datain[219:216] ^ 2);
  assign w357[24] = |(datain[215:212] ^ 12);
  assign w357[25] = |(datain[211:208] ^ 0);
  assign w357[26] = |(datain[207:204] ^ 11);
  assign w357[27] = |(datain[203:200] ^ 4);
  assign w357[28] = |(datain[199:196] ^ 4);
  assign w357[29] = |(datain[195:192] ^ 2);
  assign w357[30] = |(datain[191:188] ^ 12);
  assign w357[31] = |(datain[187:184] ^ 13);
  assign w357[32] = |(datain[183:180] ^ 2);
  assign w357[33] = |(datain[179:176] ^ 1);
  assign w357[34] = |(datain[175:172] ^ 11);
  assign w357[35] = |(datain[171:168] ^ 9);
  assign w357[36] = |(datain[167:164] ^ 0);
  assign w357[37] = |(datain[163:160] ^ 5);
  assign w357[38] = |(datain[159:156] ^ 0);
  assign w357[39] = |(datain[155:152] ^ 0);
  assign w357[40] = |(datain[151:148] ^ 11);
  assign w357[41] = |(datain[147:144] ^ 10);
  assign w357[42] = |(datain[143:140] ^ 6);
  assign w357[43] = |(datain[139:136] ^ 12);
  assign comp[357] = ~(|w357);
  wire [40-1:0] w358;
  assign w358[0] = |(datain[311:308] ^ 8);
  assign w358[1] = |(datain[307:304] ^ 14);
  assign w358[2] = |(datain[303:300] ^ 13);
  assign w358[3] = |(datain[299:296] ^ 11);
  assign w358[4] = |(datain[295:292] ^ 15);
  assign w358[5] = |(datain[291:288] ^ 15);
  assign w358[6] = |(datain[287:284] ^ 11);
  assign w358[7] = |(datain[283:280] ^ 7);
  assign w358[8] = |(datain[279:276] ^ 9);
  assign w358[9] = |(datain[275:272] ^ 0);
  assign w358[10] = |(datain[271:268] ^ 0);
  assign w358[11] = |(datain[267:264] ^ 0);
  assign w358[12] = |(datain[263:260] ^ 15);
  assign w358[13] = |(datain[259:256] ^ 15);
  assign w358[14] = |(datain[255:252] ^ 11);
  assign w358[15] = |(datain[251:248] ^ 7);
  assign w358[16] = |(datain[247:244] ^ 9);
  assign w358[17] = |(datain[243:240] ^ 2);
  assign w358[18] = |(datain[239:236] ^ 0);
  assign w358[19] = |(datain[235:232] ^ 0);
  assign w358[20] = |(datain[231:228] ^ 12);
  assign w358[21] = |(datain[227:224] ^ 7);
  assign w358[22] = |(datain[223:220] ^ 8);
  assign w358[23] = |(datain[219:216] ^ 7);
  assign w358[24] = |(datain[215:212] ^ 9);
  assign w358[25] = |(datain[211:208] ^ 0);
  assign w358[26] = |(datain[207:204] ^ 0);
  assign w358[27] = |(datain[203:200] ^ 0);
  assign w358[28] = |(datain[199:196] ^ 7);
  assign w358[29] = |(datain[195:192] ^ 2);
  assign w358[30] = |(datain[191:188] ^ 0);
  assign w358[31] = |(datain[187:184] ^ 2);
  assign w358[32] = |(datain[183:180] ^ 8);
  assign w358[33] = |(datain[179:176] ^ 12);
  assign w358[34] = |(datain[175:172] ^ 8);
  assign w358[35] = |(datain[171:168] ^ 15);
  assign w358[36] = |(datain[167:164] ^ 9);
  assign w358[37] = |(datain[163:160] ^ 2);
  assign w358[38] = |(datain[159:156] ^ 0);
  assign w358[39] = |(datain[155:152] ^ 0);
  assign comp[358] = ~(|w358);
  wire [28-1:0] w359;
  assign w359[0] = |(datain[311:308] ^ 12);
  assign w359[1] = |(datain[307:304] ^ 6);
  assign w359[2] = |(datain[303:300] ^ 7);
  assign w359[3] = |(datain[299:296] ^ 3);
  assign w359[4] = |(datain[295:292] ^ 0);
  assign w359[5] = |(datain[291:288] ^ 7);
  assign w359[6] = |(datain[287:284] ^ 2);
  assign w359[7] = |(datain[283:280] ^ 6);
  assign w359[8] = |(datain[279:276] ^ 12);
  assign w359[9] = |(datain[275:272] ^ 6);
  assign w359[10] = |(datain[271:268] ^ 0);
  assign w359[11] = |(datain[267:264] ^ 5);
  assign w359[12] = |(datain[263:260] ^ 12);
  assign w359[13] = |(datain[259:256] ^ 15);
  assign w359[14] = |(datain[255:252] ^ 4);
  assign w359[15] = |(datain[251:248] ^ 15);
  assign w359[16] = |(datain[247:244] ^ 14);
  assign w359[17] = |(datain[243:240] ^ 11);
  assign w359[18] = |(datain[239:236] ^ 15);
  assign w359[19] = |(datain[235:232] ^ 0);
  assign w359[20] = |(datain[231:228] ^ 2);
  assign w359[21] = |(datain[227:224] ^ 6);
  assign w359[22] = |(datain[223:220] ^ 15);
  assign w359[23] = |(datain[219:216] ^ 15);
  assign w359[24] = |(datain[215:212] ^ 0);
  assign w359[25] = |(datain[211:208] ^ 6);
  assign w359[26] = |(datain[207:204] ^ 0);
  assign w359[27] = |(datain[203:200] ^ 3);
  assign comp[359] = ~(|w359);
  wire [32-1:0] w360;
  assign w360[0] = |(datain[311:308] ^ 8);
  assign w360[1] = |(datain[307:304] ^ 12);
  assign w360[2] = |(datain[303:300] ^ 13);
  assign w360[3] = |(datain[299:296] ^ 13);
  assign w360[4] = |(datain[295:292] ^ 3);
  assign w360[5] = |(datain[291:288] ^ 3);
  assign w360[6] = |(datain[287:284] ^ 13);
  assign w360[7] = |(datain[283:280] ^ 11);
  assign w360[8] = |(datain[279:276] ^ 8);
  assign w360[9] = |(datain[275:272] ^ 14);
  assign w360[10] = |(datain[271:268] ^ 13);
  assign w360[11] = |(datain[267:264] ^ 11);
  assign w360[12] = |(datain[263:260] ^ 8);
  assign w360[13] = |(datain[259:256] ^ 11);
  assign w360[14] = |(datain[255:252] ^ 0);
  assign w360[15] = |(datain[251:248] ^ 7);
  assign w360[16] = |(datain[247:244] ^ 0);
  assign w360[17] = |(datain[243:240] ^ 11);
  assign w360[18] = |(datain[239:236] ^ 4);
  assign w360[19] = |(datain[235:232] ^ 7);
  assign w360[20] = |(datain[231:228] ^ 0);
  assign w360[21] = |(datain[227:224] ^ 2);
  assign w360[22] = |(datain[223:220] ^ 7);
  assign w360[23] = |(datain[219:216] ^ 4);
  assign w360[24] = |(datain[215:212] ^ 7);
  assign w360[25] = |(datain[211:208] ^ 4);
  assign w360[26] = |(datain[207:204] ^ 8);
  assign w360[27] = |(datain[203:200] ^ 9);
  assign w360[28] = |(datain[199:196] ^ 1);
  assign w360[29] = |(datain[195:192] ^ 15);
  assign w360[30] = |(datain[191:188] ^ 8);
  assign w360[31] = |(datain[187:184] ^ 9);
  assign comp[360] = ~(|w360);
  wire [60-1:0] w361;
  assign w361[0] = |(datain[311:308] ^ 0);
  assign w361[1] = |(datain[307:304] ^ 6);
  assign w361[2] = |(datain[303:300] ^ 15);
  assign w361[3] = |(datain[299:296] ^ 9);
  assign w361[4] = |(datain[295:292] ^ 0);
  assign w361[5] = |(datain[291:288] ^ 0);
  assign w361[6] = |(datain[287:284] ^ 0);
  assign w361[7] = |(datain[283:280] ^ 1);
  assign w361[8] = |(datain[279:276] ^ 3);
  assign w361[9] = |(datain[275:272] ^ 12);
  assign w361[10] = |(datain[271:268] ^ 13);
  assign w361[11] = |(datain[267:264] ^ 3);
  assign w361[12] = |(datain[263:260] ^ 7);
  assign w361[13] = |(datain[259:256] ^ 5);
  assign w361[14] = |(datain[255:252] ^ 0);
  assign w361[15] = |(datain[251:248] ^ 6);
  assign w361[16] = |(datain[247:244] ^ 2);
  assign w361[17] = |(datain[243:240] ^ 14);
  assign w361[18] = |(datain[239:236] ^ 12);
  assign w361[19] = |(datain[235:232] ^ 6);
  assign w361[20] = |(datain[231:228] ^ 0);
  assign w361[21] = |(datain[227:224] ^ 6);
  assign w361[22] = |(datain[223:220] ^ 15);
  assign w361[23] = |(datain[219:216] ^ 9);
  assign w361[24] = |(datain[215:212] ^ 0);
  assign w361[25] = |(datain[211:208] ^ 0);
  assign w361[26] = |(datain[207:204] ^ 0);
  assign w361[27] = |(datain[203:200] ^ 0);
  assign w361[28] = |(datain[199:196] ^ 11);
  assign w361[29] = |(datain[195:192] ^ 11);
  assign w361[30] = |(datain[191:188] ^ 4);
  assign w361[31] = |(datain[187:184] ^ 0);
  assign w361[32] = |(datain[183:180] ^ 0);
  assign w361[33] = |(datain[179:176] ^ 0);
  assign w361[34] = |(datain[175:172] ^ 8);
  assign w361[35] = |(datain[171:168] ^ 14);
  assign w361[36] = |(datain[167:164] ^ 13);
  assign w361[37] = |(datain[163:160] ^ 11);
  assign w361[38] = |(datain[159:156] ^ 3);
  assign w361[39] = |(datain[155:152] ^ 3);
  assign w361[40] = |(datain[151:148] ^ 13);
  assign w361[41] = |(datain[147:144] ^ 11);
  assign w361[42] = |(datain[143:140] ^ 8);
  assign w361[43] = |(datain[139:136] ^ 10);
  assign w361[44] = |(datain[135:132] ^ 4);
  assign w361[45] = |(datain[131:128] ^ 7);
  assign w361[46] = |(datain[127:124] ^ 1);
  assign w361[47] = |(datain[123:120] ^ 7);
  assign w361[48] = |(datain[119:116] ^ 2);
  assign w361[49] = |(datain[115:112] ^ 4);
  assign w361[50] = |(datain[111:108] ^ 0);
  assign w361[51] = |(datain[107:104] ^ 12);
  assign w361[52] = |(datain[103:100] ^ 3);
  assign w361[53] = |(datain[99:96] ^ 12);
  assign w361[54] = |(datain[95:92] ^ 0);
  assign w361[55] = |(datain[91:88] ^ 12);
  assign w361[56] = |(datain[87:84] ^ 7);
  assign w361[57] = |(datain[83:80] ^ 5);
  assign w361[58] = |(datain[79:76] ^ 4);
  assign w361[59] = |(datain[75:72] ^ 1);
  assign comp[361] = ~(|w361);
  wire [32-1:0] w362;
  assign w362[0] = |(datain[311:308] ^ 14);
  assign w362[1] = |(datain[307:304] ^ 8);
  assign w362[2] = |(datain[303:300] ^ 0);
  assign w362[3] = |(datain[299:296] ^ 0);
  assign w362[4] = |(datain[295:292] ^ 0);
  assign w362[5] = |(datain[291:288] ^ 0);
  assign w362[6] = |(datain[287:284] ^ 5);
  assign w362[7] = |(datain[283:280] ^ 14);
  assign w362[8] = |(datain[279:276] ^ 8);
  assign w362[9] = |(datain[275:272] ^ 1);
  assign w362[10] = |(datain[271:268] ^ 14);
  assign w362[11] = |(datain[267:264] ^ 14);
  assign w362[12] = |(datain[263:260] ^ 2);
  assign w362[13] = |(datain[259:256] ^ 9);
  assign w362[14] = |(datain[255:252] ^ 0);
  assign w362[15] = |(datain[251:248] ^ 1);
  assign w362[16] = |(datain[247:244] ^ 11);
  assign w362[17] = |(datain[243:240] ^ 9);
  assign w362[18] = |(datain[239:236] ^ 6);
  assign w362[19] = |(datain[235:232] ^ 8);
  assign w362[20] = |(datain[231:228] ^ 0);
  assign w362[21] = |(datain[227:224] ^ 5);
  assign w362[22] = |(datain[223:220] ^ 8);
  assign w362[23] = |(datain[219:216] ^ 14);
  assign w362[24] = |(datain[215:212] ^ 12);
  assign w362[25] = |(datain[211:208] ^ 5);
  assign w362[26] = |(datain[207:204] ^ 11);
  assign w362[27] = |(datain[203:200] ^ 11);
  assign w362[28] = |(datain[199:196] ^ 15);
  assign w362[29] = |(datain[195:192] ^ 15);
  assign w362[30] = |(datain[191:188] ^ 15);
  assign w362[31] = |(datain[187:184] ^ 15);
  assign comp[362] = ~(|w362);
  wire [42-1:0] w363;
  assign w363[0] = |(datain[311:308] ^ 7);
  assign w363[1] = |(datain[307:304] ^ 4);
  assign w363[2] = |(datain[303:300] ^ 0);
  assign w363[3] = |(datain[299:296] ^ 12);
  assign w363[4] = |(datain[295:292] ^ 8);
  assign w363[5] = |(datain[291:288] ^ 0);
  assign w363[6] = |(datain[287:284] ^ 7);
  assign w363[7] = |(datain[283:280] ^ 12);
  assign w363[8] = |(datain[279:276] ^ 15);
  assign w363[9] = |(datain[275:272] ^ 14);
  assign w363[10] = |(datain[271:268] ^ 3);
  assign w363[11] = |(datain[267:264] ^ 11);
  assign w363[12] = |(datain[263:260] ^ 7);
  assign w363[13] = |(datain[259:256] ^ 4);
  assign w363[14] = |(datain[255:252] ^ 0);
  assign w363[15] = |(datain[251:248] ^ 6);
  assign w363[16] = |(datain[247:244] ^ 10);
  assign w363[17] = |(datain[243:240] ^ 10);
  assign w363[18] = |(datain[239:236] ^ 14);
  assign w363[19] = |(datain[235:232] ^ 8);
  assign w363[20] = |(datain[231:228] ^ 0);
  assign w363[21] = |(datain[227:224] ^ 3);
  assign w363[22] = |(datain[223:220] ^ 0);
  assign w363[23] = |(datain[219:216] ^ 0);
  assign w363[24] = |(datain[215:212] ^ 0);
  assign w363[25] = |(datain[211:208] ^ 14);
  assign w363[26] = |(datain[207:204] ^ 1);
  assign w363[27] = |(datain[203:200] ^ 15);
  assign w363[28] = |(datain[199:196] ^ 12);
  assign w363[29] = |(datain[195:192] ^ 3);
  assign w363[30] = |(datain[191:188] ^ 5);
  assign w363[31] = |(datain[187:184] ^ 6);
  assign w363[32] = |(datain[183:180] ^ 5);
  assign w363[33] = |(datain[179:176] ^ 1);
  assign w363[34] = |(datain[175:172] ^ 1);
  assign w363[35] = |(datain[171:168] ^ 14);
  assign w363[36] = |(datain[167:164] ^ 0);
  assign w363[37] = |(datain[163:160] ^ 6);
  assign w363[38] = |(datain[159:156] ^ 0);
  assign w363[39] = |(datain[155:152] ^ 14);
  assign w363[40] = |(datain[151:148] ^ 1);
  assign w363[41] = |(datain[147:144] ^ 15);
  assign comp[363] = ~(|w363);
  wire [28-1:0] w364;
  assign w364[0] = |(datain[311:308] ^ 10);
  assign w364[1] = |(datain[307:304] ^ 3);
  assign w364[2] = |(datain[303:300] ^ 0);
  assign w364[3] = |(datain[299:296] ^ 0);
  assign w364[4] = |(datain[295:292] ^ 0);
  assign w364[5] = |(datain[291:288] ^ 1);
  assign w364[6] = |(datain[287:284] ^ 8);
  assign w364[7] = |(datain[283:280] ^ 10);
  assign w364[8] = |(datain[279:276] ^ 4);
  assign w364[9] = |(datain[275:272] ^ 6);
  assign w364[10] = |(datain[271:268] ^ 1);
  assign w364[11] = |(datain[267:264] ^ 5);
  assign w364[12] = |(datain[263:260] ^ 10);
  assign w364[13] = |(datain[259:256] ^ 2);
  assign w364[14] = |(datain[255:252] ^ 0);
  assign w364[15] = |(datain[251:248] ^ 2);
  assign w364[16] = |(datain[247:244] ^ 0);
  assign w364[17] = |(datain[243:240] ^ 1);
  assign w364[18] = |(datain[239:236] ^ 10);
  assign w364[19] = |(datain[235:232] ^ 1);
  assign w364[20] = |(datain[231:228] ^ 2);
  assign w364[21] = |(datain[227:224] ^ 12);
  assign w364[22] = |(datain[223:220] ^ 0);
  assign w364[23] = |(datain[219:216] ^ 0);
  assign w364[24] = |(datain[215:212] ^ 8);
  assign w364[25] = |(datain[211:208] ^ 14);
  assign w364[26] = |(datain[207:204] ^ 12);
  assign w364[27] = |(datain[203:200] ^ 0);
  assign comp[364] = ~(|w364);
  wire [42-1:0] w365;
  assign w365[0] = |(datain[311:308] ^ 7);
  assign w365[1] = |(datain[307:304] ^ 4);
  assign w365[2] = |(datain[303:300] ^ 0);
  assign w365[3] = |(datain[299:296] ^ 8);
  assign w365[4] = |(datain[295:292] ^ 2);
  assign w365[5] = |(datain[291:288] ^ 6);
  assign w365[6] = |(datain[287:284] ^ 8);
  assign w365[7] = |(datain[283:280] ^ 0);
  assign w365[8] = |(datain[279:276] ^ 7);
  assign w365[9] = |(datain[275:272] ^ 13);
  assign w365[10] = |(datain[271:268] ^ 15);
  assign w365[11] = |(datain[267:264] ^ 14);
  assign w365[12] = |(datain[263:260] ^ 0);
  assign w365[13] = |(datain[259:256] ^ 0);
  assign w365[14] = |(datain[255:252] ^ 7);
  assign w365[15] = |(datain[251:248] ^ 4);
  assign w365[16] = |(datain[247:244] ^ 0);
  assign w365[17] = |(datain[243:240] ^ 5);
  assign w365[18] = |(datain[239:236] ^ 4);
  assign w365[19] = |(datain[235:232] ^ 1);
  assign w365[20] = |(datain[231:228] ^ 10);
  assign w365[21] = |(datain[227:224] ^ 10);
  assign w365[22] = |(datain[223:220] ^ 14);
  assign w365[23] = |(datain[219:216] ^ 8);
  assign w365[24] = |(datain[215:212] ^ 0);
  assign w365[25] = |(datain[211:208] ^ 15);
  assign w365[26] = |(datain[207:204] ^ 0);
  assign w365[27] = |(datain[203:200] ^ 0);
  assign w365[28] = |(datain[199:196] ^ 0);
  assign w365[29] = |(datain[195:192] ^ 14);
  assign w365[30] = |(datain[191:188] ^ 1);
  assign w365[31] = |(datain[187:184] ^ 15);
  assign w365[32] = |(datain[183:180] ^ 11);
  assign w365[33] = |(datain[179:176] ^ 10);
  assign w365[34] = |(datain[175:172] ^ 8);
  assign w365[35] = |(datain[171:168] ^ 0);
  assign w365[36] = |(datain[167:164] ^ 0);
  assign w365[37] = |(datain[163:160] ^ 0);
  assign w365[38] = |(datain[159:156] ^ 11);
  assign w365[39] = |(datain[155:152] ^ 4);
  assign w365[40] = |(datain[151:148] ^ 1);
  assign w365[41] = |(datain[147:144] ^ 10);
  assign comp[365] = ~(|w365);
  wire [30-1:0] w366;
  assign w366[0] = |(datain[311:308] ^ 10);
  assign w366[1] = |(datain[307:304] ^ 13);
  assign w366[2] = |(datain[303:300] ^ 0);
  assign w366[3] = |(datain[299:296] ^ 1);
  assign w366[4] = |(datain[295:292] ^ 8);
  assign w366[5] = |(datain[291:288] ^ 11);
  assign w366[6] = |(datain[287:284] ^ 13);
  assign w366[7] = |(datain[283:280] ^ 5);
  assign w366[8] = |(datain[279:276] ^ 8);
  assign w366[9] = |(datain[275:272] ^ 3);
  assign w366[10] = |(datain[271:268] ^ 14);
  assign w366[11] = |(datain[267:264] ^ 10);
  assign w366[12] = |(datain[263:260] ^ 0);
  assign w366[13] = |(datain[259:256] ^ 4);
  assign w366[14] = |(datain[255:252] ^ 11);
  assign w366[15] = |(datain[251:248] ^ 4);
  assign w366[16] = |(datain[247:244] ^ 4);
  assign w366[17] = |(datain[243:240] ^ 0);
  assign w366[18] = |(datain[239:236] ^ 12);
  assign w366[19] = |(datain[235:232] ^ 13);
  assign w366[20] = |(datain[231:228] ^ 2);
  assign w366[21] = |(datain[227:224] ^ 1);
  assign w366[22] = |(datain[223:220] ^ 3);
  assign w366[23] = |(datain[219:216] ^ 3);
  assign w366[24] = |(datain[215:212] ^ 15);
  assign w366[25] = |(datain[211:208] ^ 15);
  assign w366[26] = |(datain[207:204] ^ 14);
  assign w366[27] = |(datain[203:200] ^ 11);
  assign w366[28] = |(datain[199:196] ^ 0);
  assign w366[29] = |(datain[195:192] ^ 3);
  assign comp[366] = ~(|w366);
  wire [28-1:0] w367;
  assign w367[0] = |(datain[311:308] ^ 0);
  assign w367[1] = |(datain[307:304] ^ 1);
  assign w367[2] = |(datain[303:300] ^ 8);
  assign w367[3] = |(datain[299:296] ^ 11);
  assign w367[4] = |(datain[295:292] ^ 13);
  assign w367[5] = |(datain[291:288] ^ 5);
  assign w367[6] = |(datain[287:284] ^ 8);
  assign w367[7] = |(datain[283:280] ^ 3);
  assign w367[8] = |(datain[279:276] ^ 14);
  assign w367[9] = |(datain[275:272] ^ 10);
  assign w367[10] = |(datain[271:268] ^ 0);
  assign w367[11] = |(datain[267:264] ^ 8);
  assign w367[12] = |(datain[263:260] ^ 11);
  assign w367[13] = |(datain[259:256] ^ 4);
  assign w367[14] = |(datain[255:252] ^ 4);
  assign w367[15] = |(datain[251:248] ^ 0);
  assign w367[16] = |(datain[247:244] ^ 12);
  assign w367[17] = |(datain[243:240] ^ 13);
  assign w367[18] = |(datain[239:236] ^ 2);
  assign w367[19] = |(datain[235:232] ^ 1);
  assign w367[20] = |(datain[231:228] ^ 3);
  assign w367[21] = |(datain[227:224] ^ 3);
  assign w367[22] = |(datain[223:220] ^ 15);
  assign w367[23] = |(datain[219:216] ^ 15);
  assign w367[24] = |(datain[215:212] ^ 14);
  assign w367[25] = |(datain[211:208] ^ 11);
  assign w367[26] = |(datain[207:204] ^ 0);
  assign w367[27] = |(datain[203:200] ^ 3);
  assign comp[367] = ~(|w367);
  wire [30-1:0] w368;
  assign w368[0] = |(datain[311:308] ^ 3);
  assign w368[1] = |(datain[307:304] ^ 15);
  assign w368[2] = |(datain[303:300] ^ 0);
  assign w368[3] = |(datain[299:296] ^ 2);
  assign w368[4] = |(datain[295:292] ^ 8);
  assign w368[5] = |(datain[291:288] ^ 11);
  assign w368[6] = |(datain[287:284] ^ 13);
  assign w368[7] = |(datain[283:280] ^ 5);
  assign w368[8] = |(datain[279:276] ^ 8);
  assign w368[9] = |(datain[275:272] ^ 3);
  assign w368[10] = |(datain[271:268] ^ 14);
  assign w368[11] = |(datain[267:264] ^ 10);
  assign w368[12] = |(datain[263:260] ^ 0);
  assign w368[13] = |(datain[259:256] ^ 14);
  assign w368[14] = |(datain[255:252] ^ 11);
  assign w368[15] = |(datain[251:248] ^ 4);
  assign w368[16] = |(datain[247:244] ^ 4);
  assign w368[17] = |(datain[243:240] ^ 0);
  assign w368[18] = |(datain[239:236] ^ 12);
  assign w368[19] = |(datain[235:232] ^ 13);
  assign w368[20] = |(datain[231:228] ^ 2);
  assign w368[21] = |(datain[227:224] ^ 1);
  assign w368[22] = |(datain[223:220] ^ 3);
  assign w368[23] = |(datain[219:216] ^ 3);
  assign w368[24] = |(datain[215:212] ^ 15);
  assign w368[25] = |(datain[211:208] ^ 15);
  assign w368[26] = |(datain[207:204] ^ 14);
  assign w368[27] = |(datain[203:200] ^ 11);
  assign w368[28] = |(datain[199:196] ^ 0);
  assign w368[29] = |(datain[195:192] ^ 3);
  assign comp[368] = ~(|w368);
  wire [30-1:0] w369;
  assign w369[0] = |(datain[311:308] ^ 5);
  assign w369[1] = |(datain[307:304] ^ 14);
  assign w369[2] = |(datain[303:300] ^ 0);
  assign w369[3] = |(datain[299:296] ^ 2);
  assign w369[4] = |(datain[295:292] ^ 8);
  assign w369[5] = |(datain[291:288] ^ 11);
  assign w369[6] = |(datain[287:284] ^ 13);
  assign w369[7] = |(datain[283:280] ^ 5);
  assign w369[8] = |(datain[279:276] ^ 8);
  assign w369[9] = |(datain[275:272] ^ 3);
  assign w369[10] = |(datain[271:268] ^ 14);
  assign w369[11] = |(datain[267:264] ^ 10);
  assign w369[12] = |(datain[263:260] ^ 0);
  assign w369[13] = |(datain[259:256] ^ 8);
  assign w369[14] = |(datain[255:252] ^ 11);
  assign w369[15] = |(datain[251:248] ^ 4);
  assign w369[16] = |(datain[247:244] ^ 4);
  assign w369[17] = |(datain[243:240] ^ 0);
  assign w369[18] = |(datain[239:236] ^ 12);
  assign w369[19] = |(datain[235:232] ^ 13);
  assign w369[20] = |(datain[231:228] ^ 2);
  assign w369[21] = |(datain[227:224] ^ 1);
  assign w369[22] = |(datain[223:220] ^ 3);
  assign w369[23] = |(datain[219:216] ^ 3);
  assign w369[24] = |(datain[215:212] ^ 15);
  assign w369[25] = |(datain[211:208] ^ 15);
  assign w369[26] = |(datain[207:204] ^ 14);
  assign w369[27] = |(datain[203:200] ^ 11);
  assign w369[28] = |(datain[199:196] ^ 0);
  assign w369[29] = |(datain[195:192] ^ 3);
  assign comp[369] = ~(|w369);
  wire [38-1:0] w370;
  assign w370[0] = |(datain[311:308] ^ 15);
  assign w370[1] = |(datain[307:304] ^ 11);
  assign w370[2] = |(datain[303:300] ^ 4);
  assign w370[3] = |(datain[299:296] ^ 0);
  assign w370[4] = |(datain[295:292] ^ 2);
  assign w370[5] = |(datain[291:288] ^ 15);
  assign w370[6] = |(datain[287:284] ^ 3);
  assign w370[7] = |(datain[283:280] ^ 11);
  assign w370[8] = |(datain[279:276] ^ 12);
  assign w370[9] = |(datain[275:272] ^ 3);
  assign w370[10] = |(datain[271:268] ^ 11);
  assign w370[11] = |(datain[267:264] ^ 9);
  assign w370[12] = |(datain[263:260] ^ 0);
  assign w370[13] = |(datain[259:256] ^ 3);
  assign w370[14] = |(datain[255:252] ^ 0);
  assign w370[15] = |(datain[251:248] ^ 0);
  assign w370[16] = |(datain[247:244] ^ 5);
  assign w370[17] = |(datain[243:240] ^ 0);
  assign w370[18] = |(datain[239:236] ^ 5);
  assign w370[19] = |(datain[235:232] ^ 3);
  assign w370[20] = |(datain[231:228] ^ 5);
  assign w370[21] = |(datain[227:224] ^ 8);
  assign w370[22] = |(datain[223:220] ^ 5);
  assign w370[23] = |(datain[219:216] ^ 11);
  assign w370[24] = |(datain[215:212] ^ 9);
  assign w370[25] = |(datain[211:208] ^ 3);
  assign w370[26] = |(datain[207:204] ^ 14);
  assign w370[27] = |(datain[203:200] ^ 2);
  assign w370[28] = |(datain[199:196] ^ 15);
  assign w370[29] = |(datain[195:192] ^ 9);
  assign w370[30] = |(datain[191:188] ^ 14);
  assign w370[31] = |(datain[187:184] ^ 8);
  assign w370[32] = |(datain[183:180] ^ 0);
  assign w370[33] = |(datain[179:176] ^ 0);
  assign w370[34] = |(datain[175:172] ^ 0);
  assign w370[35] = |(datain[171:168] ^ 0);
  assign w370[36] = |(datain[167:164] ^ 11);
  assign w370[37] = |(datain[163:160] ^ 11);
  assign comp[370] = ~(|w370);
  wire [42-1:0] w371;
  assign w371[0] = |(datain[311:308] ^ 5);
  assign w371[1] = |(datain[307:304] ^ 11);
  assign w371[2] = |(datain[303:300] ^ 11);
  assign w371[3] = |(datain[299:296] ^ 4);
  assign w371[4] = |(datain[295:292] ^ 0);
  assign w371[5] = |(datain[291:288] ^ 9);
  assign w371[6] = |(datain[287:284] ^ 8);
  assign w371[7] = |(datain[283:280] ^ 0);
  assign w371[8] = |(datain[279:276] ^ 12);
  assign w371[9] = |(datain[275:272] ^ 4);
  assign w371[10] = |(datain[271:268] ^ 3);
  assign w371[11] = |(datain[267:264] ^ 7);
  assign w371[12] = |(datain[263:260] ^ 11);
  assign w371[13] = |(datain[259:256] ^ 9);
  assign w371[14] = |(datain[255:252] ^ 7);
  assign w371[15] = |(datain[251:248] ^ 7);
  assign w371[16] = |(datain[247:244] ^ 0);
  assign w371[17] = |(datain[243:240] ^ 7);
  assign w371[18] = |(datain[239:236] ^ 8);
  assign w371[19] = |(datain[235:232] ^ 13);
  assign w371[20] = |(datain[231:228] ^ 9);
  assign w371[21] = |(datain[227:224] ^ 6);
  assign w371[22] = |(datain[223:220] ^ 0);
  assign w371[23] = |(datain[219:216] ^ 11);
  assign w371[24] = |(datain[215:212] ^ 0);
  assign w371[25] = |(datain[211:208] ^ 1);
  assign w371[26] = |(datain[207:204] ^ 12);
  assign w371[27] = |(datain[203:200] ^ 13);
  assign w371[28] = |(datain[199:196] ^ 2);
  assign w371[29] = |(datain[195:192] ^ 1);
  assign w371[30] = |(datain[191:188] ^ 14);
  assign w371[31] = |(datain[187:184] ^ 8);
  assign w371[32] = |(datain[183:180] ^ 0);
  assign w371[33] = |(datain[179:176] ^ 5);
  assign w371[34] = |(datain[175:172] ^ 0);
  assign w371[35] = |(datain[171:168] ^ 0);
  assign w371[36] = |(datain[167:164] ^ 14);
  assign w371[37] = |(datain[163:160] ^ 9);
  assign w371[38] = |(datain[159:156] ^ 1);
  assign w371[39] = |(datain[155:152] ^ 14);
  assign w371[40] = |(datain[151:148] ^ 15);
  assign w371[41] = |(datain[147:144] ^ 9);
  assign comp[371] = ~(|w371);
  wire [46-1:0] w372;
  assign w372[0] = |(datain[311:308] ^ 15);
  assign w372[1] = |(datain[307:304] ^ 4);
  assign w372[2] = |(datain[303:300] ^ 8);
  assign w372[3] = |(datain[299:296] ^ 11);
  assign w372[4] = |(datain[295:292] ^ 7);
  assign w372[5] = |(datain[291:288] ^ 4);
  assign w372[6] = |(datain[287:284] ^ 15);
  assign w372[7] = |(datain[283:280] ^ 14);
  assign w372[8] = |(datain[279:276] ^ 8);
  assign w372[9] = |(datain[275:272] ^ 1);
  assign w372[10] = |(datain[271:268] ^ 14);
  assign w372[11] = |(datain[267:264] ^ 14);
  assign w372[12] = |(datain[263:260] ^ 0);
  assign w372[13] = |(datain[259:256] ^ 4);
  assign w372[14] = |(datain[255:252] ^ 0);
  assign w372[15] = |(datain[251:248] ^ 1);
  assign w372[16] = |(datain[247:244] ^ 1);
  assign w372[17] = |(datain[243:240] ^ 14);
  assign w372[18] = |(datain[239:236] ^ 0);
  assign w372[19] = |(datain[235:232] ^ 6);
  assign w372[20] = |(datain[231:228] ^ 5);
  assign w372[21] = |(datain[227:224] ^ 0);
  assign w372[22] = |(datain[223:220] ^ 8);
  assign w372[23] = |(datain[219:216] ^ 11);
  assign w372[24] = |(datain[215:212] ^ 8);
  assign w372[25] = |(datain[211:208] ^ 4);
  assign w372[26] = |(datain[207:204] ^ 6);
  assign w372[27] = |(datain[203:200] ^ 12);
  assign w372[28] = |(datain[199:196] ^ 0);
  assign w372[29] = |(datain[195:192] ^ 2);
  assign w372[30] = |(datain[191:188] ^ 10);
  assign w372[31] = |(datain[187:184] ^ 3);
  assign w372[32] = |(datain[183:180] ^ 0);
  assign w372[33] = |(datain[179:176] ^ 0);
  assign w372[34] = |(datain[175:172] ^ 0);
  assign w372[35] = |(datain[171:168] ^ 1);
  assign w372[36] = |(datain[167:164] ^ 8);
  assign w372[37] = |(datain[163:160] ^ 11);
  assign w372[38] = |(datain[159:156] ^ 8);
  assign w372[39] = |(datain[155:152] ^ 4);
  assign w372[40] = |(datain[151:148] ^ 6);
  assign w372[41] = |(datain[147:144] ^ 14);
  assign w372[42] = |(datain[143:140] ^ 0);
  assign w372[43] = |(datain[139:136] ^ 2);
  assign w372[44] = |(datain[135:132] ^ 10);
  assign w372[45] = |(datain[131:128] ^ 3);
  assign comp[372] = ~(|w372);
  wire [48-1:0] w373;
  assign w373[0] = |(datain[311:308] ^ 11);
  assign w373[1] = |(datain[307:304] ^ 15);
  assign w373[2] = |(datain[303:300] ^ 0);
  assign w373[3] = |(datain[299:296] ^ 0);
  assign w373[4] = |(datain[295:292] ^ 0);
  assign w373[5] = |(datain[291:288] ^ 1);
  assign w373[6] = |(datain[287:284] ^ 8);
  assign w373[7] = |(datain[283:280] ^ 13);
  assign w373[8] = |(datain[279:276] ^ 11);
  assign w373[9] = |(datain[275:272] ^ 6);
  assign w373[10] = |(datain[271:268] ^ 4);
  assign w373[11] = |(datain[267:264] ^ 10);
  assign w373[12] = |(datain[263:260] ^ 0);
  assign w373[13] = |(datain[259:256] ^ 3);
  assign w373[14] = |(datain[255:252] ^ 11);
  assign w373[15] = |(datain[251:248] ^ 9);
  assign w373[16] = |(datain[247:244] ^ 0);
  assign w373[17] = |(datain[243:240] ^ 3);
  assign w373[18] = |(datain[239:236] ^ 0);
  assign w373[19] = |(datain[235:232] ^ 0);
  assign w373[20] = |(datain[231:228] ^ 15);
  assign w373[21] = |(datain[227:224] ^ 3);
  assign w373[22] = |(datain[223:220] ^ 10);
  assign w373[23] = |(datain[219:216] ^ 4);
  assign w373[24] = |(datain[215:212] ^ 12);
  assign w373[25] = |(datain[211:208] ^ 6);
  assign w373[26] = |(datain[207:204] ^ 8);
  assign w373[27] = |(datain[203:200] ^ 6);
  assign w373[28] = |(datain[199:196] ^ 5);
  assign w373[29] = |(datain[195:192] ^ 10);
  assign w373[30] = |(datain[191:188] ^ 0);
  assign w373[31] = |(datain[187:184] ^ 3);
  assign w373[32] = |(datain[183:180] ^ 0);
  assign w373[33] = |(datain[179:176] ^ 0);
  assign w373[34] = |(datain[175:172] ^ 12);
  assign w373[35] = |(datain[171:168] ^ 6);
  assign w373[36] = |(datain[167:164] ^ 8);
  assign w373[37] = |(datain[163:160] ^ 6);
  assign w373[38] = |(datain[159:156] ^ 5);
  assign w373[39] = |(datain[155:152] ^ 11);
  assign w373[40] = |(datain[151:148] ^ 0);
  assign w373[41] = |(datain[147:144] ^ 3);
  assign w373[42] = |(datain[143:140] ^ 0);
  assign w373[43] = |(datain[139:136] ^ 0);
  assign w373[44] = |(datain[135:132] ^ 14);
  assign w373[45] = |(datain[131:128] ^ 8);
  assign w373[46] = |(datain[127:124] ^ 0);
  assign w373[47] = |(datain[123:120] ^ 11);
  assign comp[373] = ~(|w373);
  wire [76-1:0] w374;
  assign w374[0] = |(datain[311:308] ^ 7);
  assign w374[1] = |(datain[307:304] ^ 12);
  assign w374[2] = |(datain[303:300] ^ 8);
  assign w374[3] = |(datain[299:296] ^ 14);
  assign w374[4] = |(datain[295:292] ^ 13);
  assign w374[5] = |(datain[291:288] ^ 8);
  assign w374[6] = |(datain[287:284] ^ 10);
  assign w374[7] = |(datain[283:280] ^ 1);
  assign w374[8] = |(datain[279:276] ^ 1);
  assign w374[9] = |(datain[275:272] ^ 3);
  assign w374[10] = |(datain[271:268] ^ 0);
  assign w374[11] = |(datain[267:264] ^ 4);
  assign w374[12] = |(datain[263:260] ^ 2);
  assign w374[13] = |(datain[259:256] ^ 13);
  assign w374[14] = |(datain[255:252] ^ 0);
  assign w374[15] = |(datain[251:248] ^ 3);
  assign w374[16] = |(datain[247:244] ^ 0);
  assign w374[17] = |(datain[243:240] ^ 0);
  assign w374[18] = |(datain[239:236] ^ 10);
  assign w374[19] = |(datain[235:232] ^ 3);
  assign w374[20] = |(datain[231:228] ^ 1);
  assign w374[21] = |(datain[227:224] ^ 3);
  assign w374[22] = |(datain[223:220] ^ 0);
  assign w374[23] = |(datain[219:216] ^ 4);
  assign w374[24] = |(datain[215:212] ^ 11);
  assign w374[25] = |(datain[211:208] ^ 1);
  assign w374[26] = |(datain[207:204] ^ 0);
  assign w374[27] = |(datain[203:200] ^ 6);
  assign w374[28] = |(datain[199:196] ^ 13);
  assign w374[29] = |(datain[195:192] ^ 3);
  assign w374[30] = |(datain[191:188] ^ 14);
  assign w374[31] = |(datain[187:184] ^ 0);
  assign w374[32] = |(datain[183:180] ^ 8);
  assign w374[33] = |(datain[179:176] ^ 14);
  assign w374[34] = |(datain[175:172] ^ 12);
  assign w374[35] = |(datain[171:168] ^ 0);
  assign w374[36] = |(datain[167:164] ^ 11);
  assign w374[37] = |(datain[163:160] ^ 14);
  assign w374[38] = |(datain[159:156] ^ 0);
  assign w374[39] = |(datain[155:152] ^ 0);
  assign w374[40] = |(datain[151:148] ^ 7);
  assign w374[41] = |(datain[147:144] ^ 12);
  assign w374[42] = |(datain[143:140] ^ 11);
  assign w374[43] = |(datain[139:136] ^ 15);
  assign w374[44] = |(datain[135:132] ^ 0);
  assign w374[45] = |(datain[131:128] ^ 0);
  assign w374[46] = |(datain[127:124] ^ 0);
  assign w374[47] = |(datain[123:120] ^ 0);
  assign w374[48] = |(datain[119:116] ^ 11);
  assign w374[49] = |(datain[115:112] ^ 9);
  assign w374[50] = |(datain[111:108] ^ 0);
  assign w374[51] = |(datain[107:104] ^ 0);
  assign w374[52] = |(datain[103:100] ^ 0);
  assign w374[53] = |(datain[99:96] ^ 1);
  assign w374[54] = |(datain[95:92] ^ 15);
  assign w374[55] = |(datain[91:88] ^ 3);
  assign w374[56] = |(datain[87:84] ^ 10);
  assign w374[57] = |(datain[83:80] ^ 5);
  assign w374[58] = |(datain[79:76] ^ 0);
  assign w374[59] = |(datain[75:72] ^ 6);
  assign w374[60] = |(datain[71:68] ^ 11);
  assign w374[61] = |(datain[67:64] ^ 8);
  assign w374[62] = |(datain[63:60] ^ 10);
  assign w374[63] = |(datain[59:56] ^ 4);
  assign w374[64] = |(datain[55:52] ^ 0);
  assign w374[65] = |(datain[51:48] ^ 0);
  assign w374[66] = |(datain[47:44] ^ 5);
  assign w374[67] = |(datain[43:40] ^ 0);
  assign w374[68] = |(datain[39:36] ^ 12);
  assign w374[69] = |(datain[35:32] ^ 11);
  assign w374[70] = |(datain[31:28] ^ 0);
  assign w374[71] = |(datain[27:24] ^ 14);
  assign w374[72] = |(datain[23:20] ^ 1);
  assign w374[73] = |(datain[19:16] ^ 15);
  assign w374[74] = |(datain[15:12] ^ 8);
  assign w374[75] = |(datain[11:8] ^ 0);
  assign comp[374] = ~(|w374);
  wire [42-1:0] w375;
  assign w375[0] = |(datain[311:308] ^ 14);
  assign w375[1] = |(datain[307:304] ^ 2);
  assign w375[2] = |(datain[303:300] ^ 1);
  assign w375[3] = |(datain[299:296] ^ 15);
  assign w375[4] = |(datain[295:292] ^ 12);
  assign w375[5] = |(datain[291:288] ^ 12);
  assign w375[6] = |(datain[287:284] ^ 4);
  assign w375[7] = |(datain[283:280] ^ 0);
  assign w375[8] = |(datain[279:276] ^ 12);
  assign w375[9] = |(datain[275:272] ^ 3);
  assign w375[10] = |(datain[271:268] ^ 15);
  assign w375[11] = |(datain[267:264] ^ 12);
  assign w375[12] = |(datain[263:260] ^ 1);
  assign w375[13] = |(datain[259:256] ^ 14);
  assign w375[14] = |(datain[255:252] ^ 0);
  assign w375[15] = |(datain[251:248] ^ 6);
  assign w375[16] = |(datain[247:244] ^ 11);
  assign w375[17] = |(datain[243:240] ^ 4);
  assign w375[18] = |(datain[239:236] ^ 5);
  assign w375[19] = |(datain[235:232] ^ 2);
  assign w375[20] = |(datain[231:228] ^ 12);
  assign w375[21] = |(datain[227:224] ^ 13);
  assign w375[22] = |(datain[223:220] ^ 2);
  assign w375[23] = |(datain[219:216] ^ 1);
  assign w375[24] = |(datain[215:212] ^ 3);
  assign w375[25] = |(datain[211:208] ^ 3);
  assign w375[26] = |(datain[207:204] ^ 14);
  assign w375[27] = |(datain[203:200] ^ 13);
  assign w375[28] = |(datain[199:196] ^ 2);
  assign w375[29] = |(datain[195:192] ^ 6);
  assign w375[30] = |(datain[191:188] ^ 8);
  assign w375[31] = |(datain[187:184] ^ 11);
  assign w375[32] = |(datain[183:180] ^ 5);
  assign w375[33] = |(datain[179:176] ^ 7);
  assign w375[34] = |(datain[175:172] ^ 15);
  assign w375[35] = |(datain[171:168] ^ 14);
  assign w375[36] = |(datain[167:164] ^ 8);
  assign w375[37] = |(datain[163:160] ^ 14);
  assign w375[38] = |(datain[159:156] ^ 13);
  assign w375[39] = |(datain[155:152] ^ 10);
  assign w375[40] = |(datain[151:148] ^ 8);
  assign w375[41] = |(datain[147:144] ^ 0);
  assign comp[375] = ~(|w375);
  wire [42-1:0] w376;
  assign w376[0] = |(datain[311:308] ^ 11);
  assign w376[1] = |(datain[307:304] ^ 4);
  assign w376[2] = |(datain[303:300] ^ 3);
  assign w376[3] = |(datain[299:296] ^ 6);
  assign w376[4] = |(datain[295:292] ^ 12);
  assign w376[5] = |(datain[291:288] ^ 12);
  assign w376[6] = |(datain[287:284] ^ 4);
  assign w376[7] = |(datain[283:280] ^ 0);
  assign w376[8] = |(datain[279:276] ^ 12);
  assign w376[9] = |(datain[275:272] ^ 3);
  assign w376[10] = |(datain[271:268] ^ 15);
  assign w376[11] = |(datain[267:264] ^ 12);
  assign w376[12] = |(datain[263:260] ^ 1);
  assign w376[13] = |(datain[259:256] ^ 14);
  assign w376[14] = |(datain[255:252] ^ 0);
  assign w376[15] = |(datain[251:248] ^ 6);
  assign w376[16] = |(datain[247:244] ^ 11);
  assign w376[17] = |(datain[243:240] ^ 4);
  assign w376[18] = |(datain[239:236] ^ 5);
  assign w376[19] = |(datain[235:232] ^ 2);
  assign w376[20] = |(datain[231:228] ^ 12);
  assign w376[21] = |(datain[227:224] ^ 13);
  assign w376[22] = |(datain[223:220] ^ 2);
  assign w376[23] = |(datain[219:216] ^ 1);
  assign w376[24] = |(datain[215:212] ^ 2);
  assign w376[25] = |(datain[211:208] ^ 6);
  assign w376[26] = |(datain[207:204] ^ 8);
  assign w376[27] = |(datain[203:200] ^ 11);
  assign w376[28] = |(datain[199:196] ^ 5);
  assign w376[29] = |(datain[195:192] ^ 7);
  assign w376[30] = |(datain[191:188] ^ 15);
  assign w376[31] = |(datain[187:184] ^ 14);
  assign w376[32] = |(datain[183:180] ^ 2);
  assign w376[33] = |(datain[179:176] ^ 14);
  assign w376[34] = |(datain[175:172] ^ 8);
  assign w376[35] = |(datain[171:168] ^ 9);
  assign w376[36] = |(datain[167:164] ^ 1);
  assign w376[37] = |(datain[163:160] ^ 6);
  assign w376[38] = |(datain[159:156] ^ 1);
  assign w376[39] = |(datain[155:152] ^ 2);
  assign w376[40] = |(datain[151:148] ^ 0);
  assign w376[41] = |(datain[147:144] ^ 5);
  assign comp[376] = ~(|w376);
  wire [44-1:0] w377;
  assign w377[0] = |(datain[311:308] ^ 11);
  assign w377[1] = |(datain[307:304] ^ 9);
  assign w377[2] = |(datain[303:300] ^ 5);
  assign w377[3] = |(datain[299:296] ^ 4);
  assign w377[4] = |(datain[295:292] ^ 0);
  assign w377[5] = |(datain[291:288] ^ 5);
  assign w377[6] = |(datain[287:284] ^ 9);
  assign w377[7] = |(datain[283:280] ^ 0);
  assign w377[8] = |(datain[279:276] ^ 8);
  assign w377[9] = |(datain[275:272] ^ 13);
  assign w377[10] = |(datain[271:268] ^ 3);
  assign w377[11] = |(datain[267:264] ^ 14);
  assign w377[12] = |(datain[263:260] ^ 2);
  assign w377[13] = |(datain[259:256] ^ 4);
  assign w377[14] = |(datain[255:252] ^ 0);
  assign w377[15] = |(datain[251:248] ^ 1);
  assign w377[16] = |(datain[247:244] ^ 2);
  assign w377[17] = |(datain[243:240] ^ 14);
  assign w377[18] = |(datain[239:236] ^ 8);
  assign w377[19] = |(datain[235:232] ^ 11);
  assign w377[20] = |(datain[231:228] ^ 3);
  assign w377[21] = |(datain[227:224] ^ 6);
  assign w377[22] = |(datain[223:220] ^ 0);
  assign w377[23] = |(datain[219:216] ^ 2);
  assign w377[24] = |(datain[215:212] ^ 0);
  assign w377[25] = |(datain[211:208] ^ 1);
  assign w377[26] = |(datain[207:204] ^ 2);
  assign w377[27] = |(datain[203:200] ^ 14);
  assign w377[28] = |(datain[199:196] ^ 3);
  assign w377[29] = |(datain[195:192] ^ 1);
  assign w377[30] = |(datain[191:188] ^ 3);
  assign w377[31] = |(datain[187:184] ^ 13);
  assign w377[32] = |(datain[183:180] ^ 2);
  assign w377[33] = |(datain[179:176] ^ 14);
  assign w377[34] = |(datain[175:172] ^ 3);
  assign w377[35] = |(datain[171:168] ^ 1);
  assign w377[36] = |(datain[167:164] ^ 3);
  assign w377[37] = |(datain[163:160] ^ 5);
  assign w377[38] = |(datain[159:156] ^ 4);
  assign w377[39] = |(datain[155:152] ^ 7);
  assign w377[40] = |(datain[151:148] ^ 14);
  assign w377[41] = |(datain[147:144] ^ 2);
  assign w377[42] = |(datain[143:140] ^ 15);
  assign w377[43] = |(datain[139:136] ^ 7);
  assign comp[377] = ~(|w377);
  wire [46-1:0] w378;
  assign w378[0] = |(datain[311:308] ^ 2);
  assign w378[1] = |(datain[307:304] ^ 4);
  assign w378[2] = |(datain[303:300] ^ 2);
  assign w378[3] = |(datain[299:296] ^ 6);
  assign w378[4] = |(datain[295:292] ^ 8);
  assign w378[5] = |(datain[291:288] ^ 8);
  assign w378[6] = |(datain[287:284] ^ 2);
  assign w378[7] = |(datain[283:280] ^ 5);
  assign w378[8] = |(datain[279:276] ^ 15);
  assign w378[9] = |(datain[275:272] ^ 3);
  assign w378[10] = |(datain[271:268] ^ 10);
  assign w378[11] = |(datain[267:264] ^ 4);
  assign w378[12] = |(datain[263:260] ^ 0);
  assign w378[13] = |(datain[259:256] ^ 6);
  assign w378[14] = |(datain[255:252] ^ 1);
  assign w378[15] = |(datain[251:248] ^ 15);
  assign w378[16] = |(datain[247:244] ^ 3);
  assign w378[17] = |(datain[243:240] ^ 3);
  assign w378[18] = |(datain[239:236] ^ 13);
  assign w378[19] = |(datain[235:232] ^ 2);
  assign w378[20] = |(datain[231:228] ^ 11);
  assign w378[21] = |(datain[227:224] ^ 8);
  assign w378[22] = |(datain[223:220] ^ 0);
  assign w378[23] = |(datain[219:216] ^ 9);
  assign w378[24] = |(datain[215:212] ^ 2);
  assign w378[25] = |(datain[211:208] ^ 5);
  assign w378[26] = |(datain[207:204] ^ 12);
  assign w378[27] = |(datain[203:200] ^ 13);
  assign w378[28] = |(datain[199:196] ^ 2);
  assign w378[29] = |(datain[195:192] ^ 1);
  assign w378[30] = |(datain[191:188] ^ 12);
  assign w378[31] = |(datain[187:184] ^ 3);
  assign w378[32] = |(datain[183:180] ^ 5);
  assign w378[33] = |(datain[179:176] ^ 0);
  assign w378[34] = |(datain[175:172] ^ 1);
  assign w378[35] = |(datain[171:168] ^ 14);
  assign w378[36] = |(datain[167:164] ^ 3);
  assign w378[37] = |(datain[163:160] ^ 3);
  assign w378[38] = |(datain[159:156] ^ 12);
  assign w378[39] = |(datain[155:152] ^ 0);
  assign w378[40] = |(datain[151:148] ^ 8);
  assign w378[41] = |(datain[147:144] ^ 14);
  assign w378[42] = |(datain[143:140] ^ 13);
  assign w378[43] = |(datain[139:136] ^ 8);
  assign w378[44] = |(datain[135:132] ^ 15);
  assign w378[45] = |(datain[131:128] ^ 6);
  assign comp[378] = ~(|w378);
  wire [74-1:0] w379;
  assign w379[0] = |(datain[311:308] ^ 12);
  assign w379[1] = |(datain[307:304] ^ 13);
  assign w379[2] = |(datain[303:300] ^ 2);
  assign w379[3] = |(datain[299:296] ^ 1);
  assign w379[4] = |(datain[295:292] ^ 11);
  assign w379[5] = |(datain[291:288] ^ 4);
  assign w379[6] = |(datain[287:284] ^ 3);
  assign w379[7] = |(datain[283:280] ^ 14);
  assign w379[8] = |(datain[279:276] ^ 12);
  assign w379[9] = |(datain[275:272] ^ 13);
  assign w379[10] = |(datain[271:268] ^ 2);
  assign w379[11] = |(datain[267:264] ^ 1);
  assign w379[12] = |(datain[263:260] ^ 5);
  assign w379[13] = |(datain[259:256] ^ 10);
  assign w379[14] = |(datain[255:252] ^ 8);
  assign w379[15] = |(datain[251:248] ^ 11);
  assign w379[16] = |(datain[247:244] ^ 13);
  assign w379[17] = |(datain[243:240] ^ 10);
  assign w379[18] = |(datain[239:236] ^ 8);
  assign w379[19] = |(datain[235:232] ^ 0);
  assign w379[20] = |(datain[231:228] ^ 7);
  assign w379[21] = |(datain[227:224] ^ 15);
  assign w379[22] = |(datain[223:220] ^ 2);
  assign w379[23] = |(datain[219:216] ^ 6);
  assign w379[24] = |(datain[215:212] ^ 0);
  assign w379[25] = |(datain[211:208] ^ 0);
  assign w379[26] = |(datain[207:204] ^ 7);
  assign w379[27] = |(datain[203:200] ^ 5);
  assign w379[28] = |(datain[199:196] ^ 0);
  assign w379[29] = |(datain[195:192] ^ 2);
  assign w379[30] = |(datain[191:188] ^ 14);
  assign w379[31] = |(datain[187:184] ^ 11);
  assign w379[32] = |(datain[183:180] ^ 0);
  assign w379[33] = |(datain[179:176] ^ 6);
  assign w379[34] = |(datain[175:172] ^ 1);
  assign w379[35] = |(datain[171:168] ^ 15);
  assign w379[36] = |(datain[167:164] ^ 11);
  assign w379[37] = |(datain[163:160] ^ 8);
  assign w379[38] = |(datain[159:156] ^ 0);
  assign w379[39] = |(datain[155:152] ^ 0);
  assign w379[40] = |(datain[151:148] ^ 0);
  assign w379[41] = |(datain[147:144] ^ 1);
  assign w379[42] = |(datain[143:140] ^ 5);
  assign w379[43] = |(datain[139:136] ^ 0);
  assign w379[44] = |(datain[135:132] ^ 12);
  assign w379[45] = |(datain[131:128] ^ 3);
  assign w379[46] = |(datain[127:124] ^ 11);
  assign w379[47] = |(datain[123:120] ^ 4);
  assign w379[48] = |(datain[119:116] ^ 0);
  assign w379[49] = |(datain[115:112] ^ 0);
  assign w379[50] = |(datain[111:108] ^ 12);
  assign w379[51] = |(datain[107:104] ^ 13);
  assign w379[52] = |(datain[103:100] ^ 1);
  assign w379[53] = |(datain[99:96] ^ 3);
  assign w379[54] = |(datain[95:92] ^ 11);
  assign w379[55] = |(datain[91:88] ^ 8);
  assign w379[56] = |(datain[87:84] ^ 0);
  assign w379[57] = |(datain[83:80] ^ 9);
  assign w379[58] = |(datain[79:76] ^ 0);
  assign w379[59] = |(datain[75:72] ^ 5);
  assign w379[60] = |(datain[71:68] ^ 11);
  assign w379[61] = |(datain[67:64] ^ 5);
  assign w379[62] = |(datain[63:60] ^ 0);
  assign w379[63] = |(datain[59:56] ^ 0);
  assign w379[64] = |(datain[55:52] ^ 11);
  assign w379[65] = |(datain[51:48] ^ 10);
  assign w379[66] = |(datain[47:44] ^ 8);
  assign w379[67] = |(datain[43:40] ^ 0);
  assign w379[68] = |(datain[39:36] ^ 0);
  assign w379[69] = |(datain[35:32] ^ 0);
  assign w379[70] = |(datain[31:28] ^ 12);
  assign w379[71] = |(datain[27:24] ^ 13);
  assign w379[72] = |(datain[23:20] ^ 1);
  assign w379[73] = |(datain[19:16] ^ 3);
  assign comp[379] = ~(|w379);
  wire [76-1:0] w380;
  assign w380[0] = |(datain[311:308] ^ 5);
  assign w380[1] = |(datain[307:304] ^ 10);
  assign w380[2] = |(datain[303:300] ^ 0);
  assign w380[3] = |(datain[299:296] ^ 0);
  assign w380[4] = |(datain[295:292] ^ 3);
  assign w380[5] = |(datain[291:288] ^ 13);
  assign w380[6] = |(datain[287:284] ^ 11);
  assign w380[7] = |(datain[283:280] ^ 0);
  assign w380[8] = |(datain[279:276] ^ 15);
  assign w380[9] = |(datain[275:272] ^ 14);
  assign w380[10] = |(datain[271:268] ^ 7);
  assign w380[11] = |(datain[267:264] ^ 7);
  assign w380[12] = |(datain[263:260] ^ 1);
  assign w380[13] = |(datain[259:256] ^ 6);
  assign w380[14] = |(datain[255:252] ^ 11);
  assign w380[15] = |(datain[251:248] ^ 4);
  assign w380[16] = |(datain[247:244] ^ 4);
  assign w380[17] = |(datain[243:240] ^ 0);
  assign w380[18] = |(datain[239:236] ^ 11);
  assign w380[19] = |(datain[235:232] ^ 9);
  assign w380[20] = |(datain[231:228] ^ 0);
  assign w380[21] = |(datain[227:224] ^ 3);
  assign w380[22] = |(datain[223:220] ^ 0);
  assign w380[23] = |(datain[219:216] ^ 1);
  assign w380[24] = |(datain[215:212] ^ 12);
  assign w380[25] = |(datain[211:208] ^ 13);
  assign w380[26] = |(datain[207:204] ^ 2);
  assign w380[27] = |(datain[203:200] ^ 1);
  assign w380[28] = |(datain[199:196] ^ 3);
  assign w380[29] = |(datain[195:192] ^ 3);
  assign w380[30] = |(datain[191:188] ^ 12);
  assign w380[31] = |(datain[187:184] ^ 9);
  assign w380[32] = |(datain[183:180] ^ 11);
  assign w380[33] = |(datain[179:176] ^ 8);
  assign w380[34] = |(datain[175:172] ^ 0);
  assign w380[35] = |(datain[171:168] ^ 0);
  assign w380[36] = |(datain[167:164] ^ 4);
  assign w380[37] = |(datain[163:160] ^ 2);
  assign w380[38] = |(datain[159:156] ^ 12);
  assign w380[39] = |(datain[155:152] ^ 13);
  assign w380[40] = |(datain[151:148] ^ 2);
  assign w380[41] = |(datain[147:144] ^ 1);
  assign w380[42] = |(datain[143:140] ^ 11);
  assign w380[43] = |(datain[139:136] ^ 2);
  assign w380[44] = |(datain[135:132] ^ 5);
  assign w380[45] = |(datain[131:128] ^ 8);
  assign w380[46] = |(datain[127:124] ^ 11);
  assign w380[47] = |(datain[123:120] ^ 1);
  assign w380[48] = |(datain[119:116] ^ 0);
  assign w380[49] = |(datain[115:112] ^ 4);
  assign w380[50] = |(datain[111:108] ^ 11);
  assign w380[51] = |(datain[107:104] ^ 4);
  assign w380[52] = |(datain[103:100] ^ 4);
  assign w380[53] = |(datain[99:96] ^ 0);
  assign w380[54] = |(datain[95:92] ^ 12);
  assign w380[55] = |(datain[91:88] ^ 13);
  assign w380[56] = |(datain[87:84] ^ 2);
  assign w380[57] = |(datain[83:80] ^ 1);
  assign w380[58] = |(datain[79:76] ^ 5);
  assign w380[59] = |(datain[75:72] ^ 10);
  assign w380[60] = |(datain[71:68] ^ 5);
  assign w380[61] = |(datain[67:64] ^ 9);
  assign w380[62] = |(datain[63:60] ^ 11);
  assign w380[63] = |(datain[59:56] ^ 8);
  assign w380[64] = |(datain[55:52] ^ 0);
  assign w380[65] = |(datain[51:48] ^ 1);
  assign w380[66] = |(datain[47:44] ^ 5);
  assign w380[67] = |(datain[43:40] ^ 7);
  assign w380[68] = |(datain[39:36] ^ 12);
  assign w380[69] = |(datain[35:32] ^ 13);
  assign w380[70] = |(datain[31:28] ^ 2);
  assign w380[71] = |(datain[27:24] ^ 1);
  assign w380[72] = |(datain[23:20] ^ 11);
  assign w380[73] = |(datain[19:16] ^ 4);
  assign w380[74] = |(datain[15:12] ^ 3);
  assign w380[75] = |(datain[11:8] ^ 14);
  assign comp[380] = ~(|w380);
  wire [76-1:0] w381;
  assign w381[0] = |(datain[311:308] ^ 12);
  assign w381[1] = |(datain[307:304] ^ 13);
  assign w381[2] = |(datain[303:300] ^ 2);
  assign w381[3] = |(datain[299:296] ^ 1);
  assign w381[4] = |(datain[295:292] ^ 2);
  assign w381[5] = |(datain[291:288] ^ 14);
  assign w381[6] = |(datain[287:284] ^ 10);
  assign w381[7] = |(datain[283:280] ^ 3);
  assign w381[8] = |(datain[279:276] ^ 5);
  assign w381[9] = |(datain[275:272] ^ 10);
  assign w381[10] = |(datain[271:268] ^ 0);
  assign w381[11] = |(datain[267:264] ^ 0);
  assign w381[12] = |(datain[263:260] ^ 3);
  assign w381[13] = |(datain[259:256] ^ 13);
  assign w381[14] = |(datain[255:252] ^ 0);
  assign w381[15] = |(datain[251:248] ^ 10);
  assign w381[16] = |(datain[247:244] ^ 0);
  assign w381[17] = |(datain[243:240] ^ 0);
  assign w381[18] = |(datain[239:236] ^ 7);
  assign w381[19] = |(datain[235:232] ^ 2);
  assign w381[20] = |(datain[231:228] ^ 1);
  assign w381[21] = |(datain[227:224] ^ 11);
  assign w381[22] = |(datain[223:220] ^ 3);
  assign w381[23] = |(datain[219:216] ^ 13);
  assign w381[24] = |(datain[215:212] ^ 2);
  assign w381[25] = |(datain[211:208] ^ 0);
  assign w381[26] = |(datain[207:204] ^ 15);
  assign w381[27] = |(datain[203:200] ^ 13);
  assign w381[28] = |(datain[199:196] ^ 7);
  assign w381[29] = |(datain[195:192] ^ 7);
  assign w381[30] = |(datain[191:188] ^ 1);
  assign w381[31] = |(datain[187:184] ^ 6);
  assign w381[32] = |(datain[183:180] ^ 11);
  assign w381[33] = |(datain[179:176] ^ 4);
  assign w381[34] = |(datain[175:172] ^ 4);
  assign w381[35] = |(datain[171:168] ^ 0);
  assign w381[36] = |(datain[167:164] ^ 11);
  assign w381[37] = |(datain[163:160] ^ 9);
  assign w381[38] = |(datain[159:156] ^ 3);
  assign w381[39] = |(datain[155:152] ^ 0);
  assign w381[40] = |(datain[151:148] ^ 0);
  assign w381[41] = |(datain[147:144] ^ 1);
  assign w381[42] = |(datain[143:140] ^ 12);
  assign w381[43] = |(datain[139:136] ^ 13);
  assign w381[44] = |(datain[135:132] ^ 2);
  assign w381[45] = |(datain[131:128] ^ 1);
  assign w381[46] = |(datain[127:124] ^ 3);
  assign w381[47] = |(datain[123:120] ^ 3);
  assign w381[48] = |(datain[119:116] ^ 12);
  assign w381[49] = |(datain[115:112] ^ 9);
  assign w381[50] = |(datain[111:108] ^ 11);
  assign w381[51] = |(datain[107:104] ^ 8);
  assign w381[52] = |(datain[103:100] ^ 0);
  assign w381[53] = |(datain[99:96] ^ 0);
  assign w381[54] = |(datain[95:92] ^ 4);
  assign w381[55] = |(datain[91:88] ^ 2);
  assign w381[56] = |(datain[87:84] ^ 12);
  assign w381[57] = |(datain[83:80] ^ 13);
  assign w381[58] = |(datain[79:76] ^ 2);
  assign w381[59] = |(datain[75:72] ^ 1);
  assign w381[60] = |(datain[71:68] ^ 11);
  assign w381[61] = |(datain[67:64] ^ 2);
  assign w381[62] = |(datain[63:60] ^ 5);
  assign w381[63] = |(datain[59:56] ^ 8);
  assign w381[64] = |(datain[55:52] ^ 11);
  assign w381[65] = |(datain[51:48] ^ 1);
  assign w381[66] = |(datain[47:44] ^ 0);
  assign w381[67] = |(datain[43:40] ^ 4);
  assign w381[68] = |(datain[39:36] ^ 11);
  assign w381[69] = |(datain[35:32] ^ 4);
  assign w381[70] = |(datain[31:28] ^ 4);
  assign w381[71] = |(datain[27:24] ^ 0);
  assign w381[72] = |(datain[23:20] ^ 12);
  assign w381[73] = |(datain[19:16] ^ 13);
  assign w381[74] = |(datain[15:12] ^ 2);
  assign w381[75] = |(datain[11:8] ^ 1);
  assign comp[381] = ~(|w381);
  wire [74-1:0] w382;
  assign w382[0] = |(datain[311:308] ^ 15);
  assign w382[1] = |(datain[307:304] ^ 4);
  assign w382[2] = |(datain[303:300] ^ 15);
  assign w382[3] = |(datain[299:296] ^ 11);
  assign w382[4] = |(datain[295:292] ^ 7);
  assign w382[5] = |(datain[291:288] ^ 7);
  assign w382[6] = |(datain[287:284] ^ 2);
  assign w382[7] = |(datain[283:280] ^ 1);
  assign w382[8] = |(datain[279:276] ^ 2);
  assign w382[9] = |(datain[275:272] ^ 14);
  assign w382[10] = |(datain[271:268] ^ 10);
  assign w382[11] = |(datain[267:264] ^ 3);
  assign w382[12] = |(datain[263:260] ^ 3);
  assign w382[13] = |(datain[259:256] ^ 15);
  assign w382[14] = |(datain[255:252] ^ 0);
  assign w382[15] = |(datain[251:248] ^ 0);
  assign w382[16] = |(datain[247:244] ^ 0);
  assign w382[17] = |(datain[243:240] ^ 5);
  assign w382[18] = |(datain[239:236] ^ 0);
  assign w382[19] = |(datain[235:232] ^ 0);
  assign w382[20] = |(datain[231:228] ^ 0);
  assign w382[21] = |(datain[227:224] ^ 1);
  assign w382[22] = |(datain[223:220] ^ 2);
  assign w382[23] = |(datain[219:216] ^ 14);
  assign w382[24] = |(datain[215:212] ^ 10);
  assign w382[25] = |(datain[211:208] ^ 3);
  assign w382[26] = |(datain[207:204] ^ 0);
  assign w382[27] = |(datain[203:200] ^ 6);
  assign w382[28] = |(datain[199:196] ^ 0);
  assign w382[29] = |(datain[195:192] ^ 0);
  assign w382[30] = |(datain[191:188] ^ 11);
  assign w382[31] = |(datain[187:184] ^ 4);
  assign w382[32] = |(datain[183:180] ^ 4);
  assign w382[33] = |(datain[179:176] ^ 0);
  assign w382[34] = |(datain[175:172] ^ 11);
  assign w382[35] = |(datain[171:168] ^ 9);
  assign w382[36] = |(datain[167:164] ^ 7);
  assign w382[37] = |(datain[163:160] ^ 6);
  assign w382[38] = |(datain[159:156] ^ 0);
  assign w382[39] = |(datain[155:152] ^ 1);
  assign w382[40] = |(datain[151:148] ^ 12);
  assign w382[41] = |(datain[147:144] ^ 13);
  assign w382[42] = |(datain[143:140] ^ 2);
  assign w382[43] = |(datain[139:136] ^ 1);
  assign w382[44] = |(datain[135:132] ^ 3);
  assign w382[45] = |(datain[131:128] ^ 3);
  assign w382[46] = |(datain[127:124] ^ 12);
  assign w382[47] = |(datain[123:120] ^ 9);
  assign w382[48] = |(datain[119:116] ^ 11);
  assign w382[49] = |(datain[115:112] ^ 8);
  assign w382[50] = |(datain[111:108] ^ 0);
  assign w382[51] = |(datain[107:104] ^ 0);
  assign w382[52] = |(datain[103:100] ^ 4);
  assign w382[53] = |(datain[99:96] ^ 2);
  assign w382[54] = |(datain[95:92] ^ 12);
  assign w382[55] = |(datain[91:88] ^ 13);
  assign w382[56] = |(datain[87:84] ^ 2);
  assign w382[57] = |(datain[83:80] ^ 1);
  assign w382[58] = |(datain[79:76] ^ 11);
  assign w382[59] = |(datain[75:72] ^ 4);
  assign w382[60] = |(datain[71:68] ^ 4);
  assign w382[61] = |(datain[67:64] ^ 0);
  assign w382[62] = |(datain[63:60] ^ 11);
  assign w382[63] = |(datain[59:56] ^ 2);
  assign w382[64] = |(datain[55:52] ^ 3);
  assign w382[65] = |(datain[51:48] ^ 13);
  assign w382[66] = |(datain[47:44] ^ 11);
  assign w382[67] = |(datain[43:40] ^ 1);
  assign w382[68] = |(datain[39:36] ^ 0);
  assign w382[69] = |(datain[35:32] ^ 4);
  assign w382[70] = |(datain[31:28] ^ 12);
  assign w382[71] = |(datain[27:24] ^ 13);
  assign w382[72] = |(datain[23:20] ^ 2);
  assign w382[73] = |(datain[19:16] ^ 1);
  assign comp[382] = ~(|w382);
  wire [72-1:0] w383;
  assign w383[0] = |(datain[311:308] ^ 0);
  assign w383[1] = |(datain[307:304] ^ 1);
  assign w383[2] = |(datain[303:300] ^ 11);
  assign w383[3] = |(datain[299:296] ^ 4);
  assign w383[4] = |(datain[295:292] ^ 4);
  assign w383[5] = |(datain[291:288] ^ 0);
  assign w383[6] = |(datain[287:284] ^ 9);
  assign w383[7] = |(datain[283:280] ^ 12);
  assign w383[8] = |(datain[279:276] ^ 2);
  assign w383[9] = |(datain[275:272] ^ 14);
  assign w383[10] = |(datain[271:268] ^ 15);
  assign w383[11] = |(datain[267:264] ^ 15);
  assign w383[12] = |(datain[263:260] ^ 1);
  assign w383[13] = |(datain[259:256] ^ 14);
  assign w383[14] = |(datain[255:252] ^ 0);
  assign w383[15] = |(datain[251:248] ^ 3);
  assign w383[16] = |(datain[247:244] ^ 0);
  assign w383[17] = |(datain[243:240] ^ 1);
  assign w383[18] = |(datain[239:236] ^ 7);
  assign w383[19] = |(datain[235:232] ^ 3);
  assign w383[20] = |(datain[231:228] ^ 0);
  assign w383[21] = |(datain[227:224] ^ 3);
  assign w383[22] = |(datain[223:220] ^ 14);
  assign w383[23] = |(datain[219:216] ^ 11);
  assign w383[24] = |(datain[215:212] ^ 1);
  assign w383[25] = |(datain[211:208] ^ 9);
  assign w383[26] = |(datain[207:204] ^ 9);
  assign w383[27] = |(datain[203:200] ^ 0);
  assign w383[28] = |(datain[199:196] ^ 11);
  assign w383[29] = |(datain[195:192] ^ 10);
  assign w383[30] = |(datain[191:188] ^ 0);
  assign w383[31] = |(datain[187:184] ^ 0);
  assign w383[32] = |(datain[183:180] ^ 0);
  assign w383[33] = |(datain[179:176] ^ 1);
  assign w383[34] = |(datain[175:172] ^ 11);
  assign w383[35] = |(datain[171:168] ^ 9);
  assign w383[36] = |(datain[167:164] ^ 14);
  assign w383[37] = |(datain[163:160] ^ 1);
  assign w383[38] = |(datain[159:156] ^ 0);
  assign w383[39] = |(datain[155:152] ^ 3);
  assign w383[40] = |(datain[151:148] ^ 2);
  assign w383[41] = |(datain[147:144] ^ 14);
  assign w383[42] = |(datain[143:140] ^ 8);
  assign w383[43] = |(datain[139:136] ^ 11);
  assign w383[44] = |(datain[135:132] ^ 1);
  assign w383[45] = |(datain[131:128] ^ 14);
  assign w383[46] = |(datain[127:124] ^ 1);
  assign w383[47] = |(datain[123:120] ^ 8);
  assign w383[48] = |(datain[119:116] ^ 0);
  assign w383[49] = |(datain[115:112] ^ 1);
  assign w383[50] = |(datain[111:108] ^ 11);
  assign w383[51] = |(datain[107:104] ^ 4);
  assign w383[52] = |(datain[103:100] ^ 4);
  assign w383[53] = |(datain[99:96] ^ 0);
  assign w383[54] = |(datain[95:92] ^ 9);
  assign w383[55] = |(datain[91:88] ^ 12);
  assign w383[56] = |(datain[87:84] ^ 2);
  assign w383[57] = |(datain[83:80] ^ 14);
  assign w383[58] = |(datain[79:76] ^ 15);
  assign w383[59] = |(datain[75:72] ^ 15);
  assign w383[60] = |(datain[71:68] ^ 1);
  assign w383[61] = |(datain[67:64] ^ 14);
  assign w383[62] = |(datain[63:60] ^ 0);
  assign w383[63] = |(datain[59:56] ^ 3);
  assign w383[64] = |(datain[55:52] ^ 0);
  assign w383[65] = |(datain[51:48] ^ 1);
  assign w383[66] = |(datain[47:44] ^ 7);
  assign w383[67] = |(datain[43:40] ^ 3);
  assign w383[68] = |(datain[39:36] ^ 0);
  assign w383[69] = |(datain[35:32] ^ 3);
  assign w383[70] = |(datain[31:28] ^ 14);
  assign w383[71] = |(datain[27:24] ^ 11);
  assign comp[383] = ~(|w383);
  wire [76-1:0] w384;
  assign w384[0] = |(datain[311:308] ^ 7);
  assign w384[1] = |(datain[307:304] ^ 12);
  assign w384[2] = |(datain[303:300] ^ 15);
  assign w384[3] = |(datain[299:296] ^ 10);
  assign w384[4] = |(datain[295:292] ^ 8);
  assign w384[5] = |(datain[291:288] ^ 11);
  assign w384[6] = |(datain[287:284] ^ 14);
  assign w384[7] = |(datain[283:280] ^ 6);
  assign w384[8] = |(datain[279:276] ^ 8);
  assign w384[9] = |(datain[275:272] ^ 14);
  assign w384[10] = |(datain[271:268] ^ 13);
  assign w384[11] = |(datain[267:264] ^ 0);
  assign w384[12] = |(datain[263:260] ^ 15);
  assign w384[13] = |(datain[259:256] ^ 11);
  assign w384[14] = |(datain[255:252] ^ 11);
  assign w384[15] = |(datain[251:248] ^ 15);
  assign w384[16] = |(datain[247:244] ^ 1);
  assign w384[17] = |(datain[243:240] ^ 3);
  assign w384[18] = |(datain[239:236] ^ 0);
  assign w384[19] = |(datain[235:232] ^ 4);
  assign w384[20] = |(datain[231:228] ^ 8);
  assign w384[21] = |(datain[227:224] ^ 3);
  assign w384[22] = |(datain[223:220] ^ 2);
  assign w384[23] = |(datain[219:216] ^ 13);
  assign w384[24] = |(datain[215:212] ^ 0);
  assign w384[25] = |(datain[211:208] ^ 2);
  assign w384[26] = |(datain[207:204] ^ 12);
  assign w384[27] = |(datain[203:200] ^ 13);
  assign w384[28] = |(datain[199:196] ^ 1);
  assign w384[29] = |(datain[195:192] ^ 2);
  assign w384[30] = |(datain[191:188] ^ 11);
  assign w384[31] = |(datain[187:184] ^ 3);
  assign w384[32] = |(datain[183:180] ^ 0);
  assign w384[33] = |(datain[179:176] ^ 6);
  assign w384[34] = |(datain[175:172] ^ 8);
  assign w384[35] = |(datain[171:168] ^ 6);
  assign w384[36] = |(datain[167:164] ^ 13);
  assign w384[37] = |(datain[163:160] ^ 9);
  assign w384[38] = |(datain[159:156] ^ 13);
  assign w384[39] = |(datain[155:152] ^ 3);
  assign w384[40] = |(datain[151:148] ^ 14);
  assign w384[41] = |(datain[147:144] ^ 0);
  assign w384[42] = |(datain[143:140] ^ 8);
  assign w384[43] = |(datain[139:136] ^ 14);
  assign w384[44] = |(datain[135:132] ^ 12);
  assign w384[45] = |(datain[131:128] ^ 0);
  assign w384[46] = |(datain[127:124] ^ 12);
  assign w384[47] = |(datain[123:120] ^ 7);
  assign w384[48] = |(datain[119:116] ^ 0);
  assign w384[49] = |(datain[115:112] ^ 6);
  assign w384[50] = |(datain[111:108] ^ 8);
  assign w384[51] = |(datain[107:104] ^ 14);
  assign w384[52] = |(datain[103:100] ^ 0);
  assign w384[53] = |(datain[99:96] ^ 0);
  assign w384[54] = |(datain[95:92] ^ 0);
  assign w384[55] = |(datain[91:88] ^ 0);
  assign w384[56] = |(datain[87:84] ^ 0);
  assign w384[57] = |(datain[83:80] ^ 1);
  assign w384[58] = |(datain[79:76] ^ 12);
  assign w384[59] = |(datain[75:72] ^ 7);
  assign w384[60] = |(datain[71:68] ^ 0);
  assign w384[61] = |(datain[67:64] ^ 6);
  assign w384[62] = |(datain[63:60] ^ 9);
  assign w384[63] = |(datain[59:56] ^ 2);
  assign w384[64] = |(datain[55:52] ^ 0);
  assign w384[65] = |(datain[51:48] ^ 0);
  assign w384[66] = |(datain[47:44] ^ 0);
  assign w384[67] = |(datain[43:40] ^ 1);
  assign w384[68] = |(datain[39:36] ^ 0);
  assign w384[69] = |(datain[35:32] ^ 1);
  assign w384[70] = |(datain[31:28] ^ 3);
  assign w384[71] = |(datain[27:24] ^ 3);
  assign w384[72] = |(datain[23:20] ^ 12);
  assign w384[73] = |(datain[19:16] ^ 0);
  assign w384[74] = |(datain[15:12] ^ 12);
  assign w384[75] = |(datain[11:8] ^ 13);
  assign comp[384] = ~(|w384);
  wire [74-1:0] w385;
  assign w385[0] = |(datain[311:308] ^ 0);
  assign w385[1] = |(datain[307:304] ^ 1);
  assign w385[2] = |(datain[303:300] ^ 7);
  assign w385[3] = |(datain[299:296] ^ 5);
  assign w385[4] = |(datain[295:292] ^ 0);
  assign w385[5] = |(datain[291:288] ^ 5);
  assign w385[6] = |(datain[287:284] ^ 11);
  assign w385[7] = |(datain[283:280] ^ 8);
  assign w385[8] = |(datain[279:276] ^ 0);
  assign w385[9] = |(datain[275:272] ^ 1);
  assign w385[10] = |(datain[271:268] ^ 4);
  assign w385[11] = |(datain[267:264] ^ 12);
  assign w385[12] = |(datain[263:260] ^ 12);
  assign w385[13] = |(datain[259:256] ^ 13);
  assign w385[14] = |(datain[255:252] ^ 2);
  assign w385[15] = |(datain[251:248] ^ 1);
  assign w385[16] = |(datain[247:244] ^ 8);
  assign w385[17] = |(datain[243:240] ^ 9);
  assign w385[18] = |(datain[239:236] ^ 1);
  assign w385[19] = |(datain[235:232] ^ 6);
  assign w385[20] = |(datain[231:228] ^ 3);
  assign w385[21] = |(datain[227:224] ^ 7);
  assign w385[22] = |(datain[223:220] ^ 0);
  assign w385[23] = |(datain[219:216] ^ 1);
  assign w385[24] = |(datain[215:212] ^ 8);
  assign w385[25] = |(datain[211:208] ^ 9);
  assign w385[26] = |(datain[207:204] ^ 0);
  assign w385[27] = |(datain[203:200] ^ 14);
  assign w385[28] = |(datain[199:196] ^ 3);
  assign w385[29] = |(datain[195:192] ^ 9);
  assign w385[30] = |(datain[191:188] ^ 0);
  assign w385[31] = |(datain[187:184] ^ 1);
  assign w385[32] = |(datain[183:180] ^ 11);
  assign w385[33] = |(datain[179:176] ^ 10);
  assign w385[34] = |(datain[175:172] ^ 3);
  assign w385[35] = |(datain[171:168] ^ 11);
  assign w385[36] = |(datain[167:164] ^ 0);
  assign w385[37] = |(datain[163:160] ^ 1);
  assign w385[38] = |(datain[159:156] ^ 3);
  assign w385[39] = |(datain[155:152] ^ 3);
  assign w385[40] = |(datain[151:148] ^ 12);
  assign w385[41] = |(datain[147:144] ^ 9);
  assign w385[42] = |(datain[143:140] ^ 11);
  assign w385[43] = |(datain[139:136] ^ 4);
  assign w385[44] = |(datain[135:132] ^ 3);
  assign w385[45] = |(datain[131:128] ^ 12);
  assign w385[46] = |(datain[127:124] ^ 12);
  assign w385[47] = |(datain[123:120] ^ 13);
  assign w385[48] = |(datain[119:116] ^ 2);
  assign w385[49] = |(datain[115:112] ^ 1);
  assign w385[50] = |(datain[111:108] ^ 8);
  assign w385[51] = |(datain[107:104] ^ 11);
  assign w385[52] = |(datain[103:100] ^ 13);
  assign w385[53] = |(datain[99:96] ^ 8);
  assign w385[54] = |(datain[95:92] ^ 11);
  assign w385[55] = |(datain[91:88] ^ 10);
  assign w385[56] = |(datain[87:84] ^ 0);
  assign w385[57] = |(datain[83:80] ^ 0);
  assign w385[58] = |(datain[79:76] ^ 0);
  assign w385[59] = |(datain[75:72] ^ 1);
  assign w385[60] = |(datain[71:68] ^ 11);
  assign w385[61] = |(datain[67:64] ^ 9);
  assign w385[62] = |(datain[63:60] ^ 4);
  assign w385[63] = |(datain[59:56] ^ 7);
  assign w385[64] = |(datain[55:52] ^ 0);
  assign w385[65] = |(datain[51:48] ^ 0);
  assign w385[66] = |(datain[47:44] ^ 11);
  assign w385[67] = |(datain[43:40] ^ 4);
  assign w385[68] = |(datain[39:36] ^ 4);
  assign w385[69] = |(datain[35:32] ^ 0);
  assign w385[70] = |(datain[31:28] ^ 12);
  assign w385[71] = |(datain[27:24] ^ 13);
  assign w385[72] = |(datain[23:20] ^ 2);
  assign w385[73] = |(datain[19:16] ^ 1);
  assign comp[385] = ~(|w385);
  wire [72-1:0] w386;
  assign w386[0] = |(datain[311:308] ^ 11);
  assign w386[1] = |(datain[307:304] ^ 4);
  assign w386[2] = |(datain[303:300] ^ 4);
  assign w386[3] = |(datain[299:296] ^ 0);
  assign w386[4] = |(datain[295:292] ^ 11);
  assign w386[5] = |(datain[291:288] ^ 10);
  assign w386[6] = |(datain[287:284] ^ 0);
  assign w386[7] = |(datain[283:280] ^ 0);
  assign w386[8] = |(datain[279:276] ^ 0);
  assign w386[9] = |(datain[275:272] ^ 2);
  assign w386[10] = |(datain[271:268] ^ 11);
  assign w386[11] = |(datain[267:264] ^ 9);
  assign w386[12] = |(datain[263:260] ^ 15);
  assign w386[13] = |(datain[259:256] ^ 11);
  assign w386[14] = |(datain[255:252] ^ 0);
  assign w386[15] = |(datain[251:248] ^ 1);
  assign w386[16] = |(datain[247:244] ^ 9);
  assign w386[17] = |(datain[243:240] ^ 0);
  assign w386[18] = |(datain[239:236] ^ 12);
  assign w386[19] = |(datain[235:232] ^ 13);
  assign w386[20] = |(datain[231:228] ^ 3);
  assign w386[21] = |(datain[227:224] ^ 8);
  assign w386[22] = |(datain[223:220] ^ 14);
  assign w386[23] = |(datain[219:216] ^ 8);
  assign w386[24] = |(datain[215:212] ^ 2);
  assign w386[25] = |(datain[211:208] ^ 3);
  assign w386[26] = |(datain[207:204] ^ 0);
  assign w386[27] = |(datain[203:200] ^ 0);
  assign w386[28] = |(datain[199:196] ^ 5);
  assign w386[29] = |(datain[195:192] ^ 9);
  assign w386[30] = |(datain[191:188] ^ 11);
  assign w386[31] = |(datain[187:184] ^ 4);
  assign w386[32] = |(datain[183:180] ^ 4);
  assign w386[33] = |(datain[179:176] ^ 0);
  assign w386[34] = |(datain[175:172] ^ 8);
  assign w386[35] = |(datain[171:168] ^ 11);
  assign w386[36] = |(datain[167:164] ^ 13);
  assign w386[37] = |(datain[163:160] ^ 6);
  assign w386[38] = |(datain[159:156] ^ 12);
  assign w386[39] = |(datain[155:152] ^ 13);
  assign w386[40] = |(datain[151:148] ^ 3);
  assign w386[41] = |(datain[147:144] ^ 8);
  assign w386[42] = |(datain[143:140] ^ 11);
  assign w386[43] = |(datain[139:136] ^ 8);
  assign w386[44] = |(datain[135:132] ^ 0);
  assign w386[45] = |(datain[131:128] ^ 0);
  assign w386[46] = |(datain[127:124] ^ 5);
  assign w386[47] = |(datain[123:120] ^ 7);
  assign w386[48] = |(datain[119:116] ^ 12);
  assign w386[49] = |(datain[115:112] ^ 13);
  assign w386[50] = |(datain[111:108] ^ 3);
  assign w386[51] = |(datain[107:104] ^ 8);
  assign w386[52] = |(datain[103:100] ^ 4);
  assign w386[53] = |(datain[99:96] ^ 0);
  assign w386[54] = |(datain[95:92] ^ 12);
  assign w386[55] = |(datain[91:88] ^ 13);
  assign w386[56] = |(datain[87:84] ^ 3);
  assign w386[57] = |(datain[83:80] ^ 8);
  assign w386[58] = |(datain[79:76] ^ 11);
  assign w386[59] = |(datain[75:72] ^ 4);
  assign w386[60] = |(datain[71:68] ^ 3);
  assign w386[61] = |(datain[67:64] ^ 14);
  assign w386[62] = |(datain[63:60] ^ 12);
  assign w386[63] = |(datain[59:56] ^ 13);
  assign w386[64] = |(datain[55:52] ^ 3);
  assign w386[65] = |(datain[51:48] ^ 8);
  assign w386[66] = |(datain[47:44] ^ 14);
  assign w386[67] = |(datain[43:40] ^ 8);
  assign w386[68] = |(datain[39:36] ^ 1);
  assign w386[69] = |(datain[35:32] ^ 12);
  assign w386[70] = |(datain[31:28] ^ 0);
  assign w386[71] = |(datain[27:24] ^ 0);
  assign comp[386] = ~(|w386);
  wire [30-1:0] w387;
  assign w387[0] = |(datain[311:308] ^ 0);
  assign w387[1] = |(datain[307:304] ^ 1);
  assign w387[2] = |(datain[303:300] ^ 8);
  assign w387[3] = |(datain[299:296] ^ 10);
  assign w387[4] = |(datain[295:292] ^ 0);
  assign w387[5] = |(datain[291:288] ^ 7);
  assign w387[6] = |(datain[287:284] ^ 8);
  assign w387[7] = |(datain[283:280] ^ 8);
  assign w387[8] = |(datain[279:276] ^ 0);
  assign w387[9] = |(datain[275:272] ^ 5);
  assign w387[10] = |(datain[271:268] ^ 8);
  assign w387[11] = |(datain[267:264] ^ 11);
  assign w387[12] = |(datain[263:260] ^ 4);
  assign w387[13] = |(datain[259:256] ^ 7);
  assign w387[14] = |(datain[255:252] ^ 0);
  assign w387[15] = |(datain[251:248] ^ 1);
  assign w387[16] = |(datain[247:244] ^ 8);
  assign w387[17] = |(datain[243:240] ^ 9);
  assign w387[18] = |(datain[239:236] ^ 4);
  assign w387[19] = |(datain[235:232] ^ 5);
  assign w387[20] = |(datain[231:228] ^ 0);
  assign w387[21] = |(datain[227:224] ^ 1);
  assign w387[22] = |(datain[223:220] ^ 15);
  assign w387[23] = |(datain[219:216] ^ 15);
  assign w387[24] = |(datain[215:212] ^ 14);
  assign w387[25] = |(datain[211:208] ^ 7);
  assign w387[26] = |(datain[207:204] ^ 12);
  assign w387[27] = |(datain[203:200] ^ 3);
  assign w387[28] = |(datain[199:196] ^ 14);
  assign w387[29] = |(datain[195:192] ^ 8);
  assign comp[387] = ~(|w387);
  wire [46-1:0] w388;
  assign w388[0] = |(datain[311:308] ^ 0);
  assign w388[1] = |(datain[307:304] ^ 1);
  assign w388[2] = |(datain[303:300] ^ 8);
  assign w388[3] = |(datain[299:296] ^ 10);
  assign w388[4] = |(datain[295:292] ^ 0);
  assign w388[5] = |(datain[291:288] ^ 7);
  assign w388[6] = |(datain[287:284] ^ 8);
  assign w388[7] = |(datain[283:280] ^ 8);
  assign w388[8] = |(datain[279:276] ^ 0);
  assign w388[9] = |(datain[275:272] ^ 5);
  assign w388[10] = |(datain[271:268] ^ 8);
  assign w388[11] = |(datain[267:264] ^ 11);
  assign w388[12] = |(datain[263:260] ^ 4);
  assign w388[13] = |(datain[259:256] ^ 7);
  assign w388[14] = |(datain[255:252] ^ 0);
  assign w388[15] = |(datain[251:248] ^ 1);
  assign w388[16] = |(datain[247:244] ^ 8);
  assign w388[17] = |(datain[243:240] ^ 9);
  assign w388[18] = |(datain[239:236] ^ 4);
  assign w388[19] = |(datain[235:232] ^ 5);
  assign w388[20] = |(datain[231:228] ^ 0);
  assign w388[21] = |(datain[227:224] ^ 1);
  assign w388[22] = |(datain[223:220] ^ 15);
  assign w388[23] = |(datain[219:216] ^ 15);
  assign w388[24] = |(datain[215:212] ^ 14);
  assign w388[25] = |(datain[211:208] ^ 7);
  assign w388[26] = |(datain[207:204] ^ 12);
  assign w388[27] = |(datain[203:200] ^ 11);
  assign w388[28] = |(datain[199:196] ^ 14);
  assign w388[29] = |(datain[195:192] ^ 8);
  assign w388[30] = |(datain[191:188] ^ 13);
  assign w388[31] = |(datain[187:184] ^ 14);
  assign w388[32] = |(datain[183:180] ^ 0);
  assign w388[33] = |(datain[179:176] ^ 0);
  assign w388[34] = |(datain[175:172] ^ 8);
  assign w388[35] = |(datain[171:168] ^ 10);
  assign w388[36] = |(datain[167:164] ^ 8);
  assign w388[37] = |(datain[163:160] ^ 4);
  assign w388[38] = |(datain[159:156] ^ 2);
  assign w388[39] = |(datain[155:152] ^ 8);
  assign w388[40] = |(datain[151:148] ^ 0);
  assign w388[41] = |(datain[147:144] ^ 4);
  assign w388[42] = |(datain[143:140] ^ 0);
  assign w388[43] = |(datain[139:136] ^ 10);
  assign w388[44] = |(datain[135:132] ^ 12);
  assign w388[45] = |(datain[131:128] ^ 0);
  assign comp[388] = ~(|w388);
  wire [44-1:0] w389;
  assign w389[0] = |(datain[311:308] ^ 13);
  assign w389[1] = |(datain[307:304] ^ 13);
  assign w389[2] = |(datain[303:300] ^ 12);
  assign w389[3] = |(datain[299:296] ^ 13);
  assign w389[4] = |(datain[295:292] ^ 2);
  assign w389[5] = |(datain[291:288] ^ 1);
  assign w389[6] = |(datain[287:284] ^ 8);
  assign w389[7] = |(datain[283:280] ^ 0);
  assign w389[8] = |(datain[279:276] ^ 15);
  assign w389[9] = |(datain[275:272] ^ 12);
  assign w389[10] = |(datain[271:268] ^ 12);
  assign w389[11] = |(datain[267:264] ^ 12);
  assign w389[12] = |(datain[263:260] ^ 7);
  assign w389[13] = |(datain[259:256] ^ 5);
  assign w389[14] = |(datain[255:252] ^ 0);
  assign w389[15] = |(datain[251:248] ^ 7);
  assign w389[16] = |(datain[247:244] ^ 3);
  assign w389[17] = |(datain[243:240] ^ 12);
  assign w389[18] = |(datain[239:236] ^ 12);
  assign w389[19] = |(datain[235:232] ^ 0);
  assign w389[20] = |(datain[231:228] ^ 7);
  assign w389[21] = |(datain[227:224] ^ 2);
  assign w389[22] = |(datain[223:220] ^ 0);
  assign w389[23] = |(datain[219:216] ^ 3);
  assign w389[24] = |(datain[215:212] ^ 14);
  assign w389[25] = |(datain[211:208] ^ 9);
  assign w389[26] = |(datain[207:204] ^ 12);
  assign w389[27] = |(datain[203:200] ^ 14);
  assign w389[28] = |(datain[199:196] ^ 0);
  assign w389[29] = |(datain[195:192] ^ 0);
  assign w389[30] = |(datain[191:188] ^ 11);
  assign w389[31] = |(datain[187:184] ^ 8);
  assign w389[32] = |(datain[183:180] ^ 0);
  assign w389[33] = |(datain[179:176] ^ 9);
  assign w389[34] = |(datain[175:172] ^ 3);
  assign w389[35] = |(datain[171:168] ^ 5);
  assign w389[36] = |(datain[167:164] ^ 12);
  assign w389[37] = |(datain[163:160] ^ 13);
  assign w389[38] = |(datain[159:156] ^ 2);
  assign w389[39] = |(datain[155:152] ^ 1);
  assign w389[40] = |(datain[151:148] ^ 2);
  assign w389[41] = |(datain[147:144] ^ 14);
  assign w389[42] = |(datain[143:140] ^ 8);
  assign w389[43] = |(datain[139:136] ^ 9);
  assign comp[389] = ~(|w389);
  wire [32-1:0] w390;
  assign w390[0] = |(datain[311:308] ^ 1);
  assign w390[1] = |(datain[307:304] ^ 15);
  assign w390[2] = |(datain[303:300] ^ 8);
  assign w390[3] = |(datain[299:296] ^ 1);
  assign w390[4] = |(datain[295:292] ^ 14);
  assign w390[5] = |(datain[291:288] ^ 14);
  assign w390[6] = |(datain[287:284] ^ 13);
  assign w390[7] = |(datain[283:280] ^ 7);
  assign w390[8] = |(datain[279:276] ^ 0);
  assign w390[9] = |(datain[275:272] ^ 4);
  assign w390[10] = |(datain[271:268] ^ 11);
  assign w390[11] = |(datain[267:264] ^ 9);
  assign w390[12] = |(datain[263:260] ^ 4);
  assign w390[13] = |(datain[259:256] ^ 14);
  assign w390[14] = |(datain[255:252] ^ 0);
  assign w390[15] = |(datain[251:248] ^ 6);
  assign w390[16] = |(datain[247:244] ^ 4);
  assign w390[17] = |(datain[243:240] ^ 1);
  assign w390[18] = |(datain[239:236] ^ 15);
  assign w390[19] = |(datain[235:232] ^ 3);
  assign w390[20] = |(datain[231:228] ^ 10);
  assign w390[21] = |(datain[227:224] ^ 4);
  assign w390[22] = |(datain[223:220] ^ 11);
  assign w390[23] = |(datain[219:216] ^ 4);
  assign w390[24] = |(datain[215:212] ^ 6);
  assign w390[25] = |(datain[211:208] ^ 2);
  assign w390[26] = |(datain[207:204] ^ 12);
  assign w390[27] = |(datain[203:200] ^ 13);
  assign w390[28] = |(datain[199:196] ^ 2);
  assign w390[29] = |(datain[195:192] ^ 1);
  assign w390[30] = |(datain[191:188] ^ 4);
  assign w390[31] = |(datain[187:184] ^ 11);
  assign comp[390] = ~(|w390);
  wire [28-1:0] w391;
  assign w391[0] = |(datain[311:308] ^ 4);
  assign w391[1] = |(datain[307:304] ^ 0);
  assign w391[2] = |(datain[303:300] ^ 11);
  assign w391[3] = |(datain[299:296] ^ 9);
  assign w391[4] = |(datain[295:292] ^ 4);
  assign w391[5] = |(datain[291:288] ^ 14);
  assign w391[6] = |(datain[287:284] ^ 0);
  assign w391[7] = |(datain[283:280] ^ 6);
  assign w391[8] = |(datain[279:276] ^ 11);
  assign w391[9] = |(datain[275:272] ^ 10);
  assign w391[10] = |(datain[271:268] ^ 0);
  assign w391[11] = |(datain[267:264] ^ 0);
  assign w391[12] = |(datain[263:260] ^ 0);
  assign w391[13] = |(datain[259:256] ^ 1);
  assign w391[14] = |(datain[255:252] ^ 14);
  assign w391[15] = |(datain[251:248] ^ 8);
  assign w391[16] = |(datain[247:244] ^ 5);
  assign w391[17] = |(datain[243:240] ^ 10);
  assign w391[18] = |(datain[239:236] ^ 0);
  assign w391[19] = |(datain[235:232] ^ 0);
  assign w391[20] = |(datain[231:228] ^ 14);
  assign w391[21] = |(datain[227:224] ^ 11);
  assign w391[22] = |(datain[223:220] ^ 5);
  assign w391[23] = |(datain[219:216] ^ 1);
  assign w391[24] = |(datain[215:212] ^ 9);
  assign w391[25] = |(datain[211:208] ^ 0);
  assign w391[26] = |(datain[207:204] ^ 11);
  assign w391[27] = |(datain[203:200] ^ 8);
  assign comp[391] = ~(|w391);
  wire [44-1:0] w392;
  assign w392[0] = |(datain[311:308] ^ 7);
  assign w392[1] = |(datain[307:304] ^ 6);
  assign w392[2] = |(datain[303:300] ^ 15);
  assign w392[3] = |(datain[299:296] ^ 10);
  assign w392[4] = |(datain[295:292] ^ 9);
  assign w392[5] = |(datain[291:288] ^ 10);
  assign w392[6] = |(datain[287:284] ^ 0);
  assign w392[7] = |(datain[283:280] ^ 2);
  assign w392[8] = |(datain[279:276] ^ 3);
  assign w392[9] = |(datain[275:272] ^ 6);
  assign w392[10] = |(datain[271:268] ^ 8);
  assign w392[11] = |(datain[267:264] ^ 1);
  assign w392[12] = |(datain[263:260] ^ 7);
  assign w392[13] = |(datain[259:256] ^ 14);
  assign w392[14] = |(datain[255:252] ^ 15);
  assign w392[15] = |(datain[251:248] ^ 10);
  assign w392[16] = |(datain[247:244] ^ 12);
  assign w392[17] = |(datain[243:240] ^ 0);
  assign w392[18] = |(datain[239:236] ^ 4);
  assign w392[19] = |(datain[235:232] ^ 15);
  assign w392[20] = |(datain[231:228] ^ 7);
  assign w392[21] = |(datain[227:224] ^ 5);
  assign w392[22] = |(datain[223:220] ^ 0);
  assign w392[23] = |(datain[219:216] ^ 3);
  assign w392[24] = |(datain[215:212] ^ 14);
  assign w392[25] = |(datain[211:208] ^ 9);
  assign w392[26] = |(datain[207:204] ^ 1);
  assign w392[27] = |(datain[203:200] ^ 1);
  assign w392[28] = |(datain[199:196] ^ 0);
  assign w392[29] = |(datain[195:192] ^ 0);
  assign w392[30] = |(datain[191:188] ^ 3);
  assign w392[31] = |(datain[187:184] ^ 6);
  assign w392[32] = |(datain[183:180] ^ 8);
  assign w392[33] = |(datain[179:176] ^ 1);
  assign w392[34] = |(datain[175:172] ^ 7);
  assign w392[35] = |(datain[171:168] ^ 14);
  assign w392[36] = |(datain[167:164] ^ 15);
  assign w392[37] = |(datain[163:160] ^ 10);
  assign w392[38] = |(datain[159:156] ^ 13);
  assign w392[39] = |(datain[155:152] ^ 7);
  assign w392[40] = |(datain[151:148] ^ 5);
  assign w392[41] = |(datain[147:144] ^ 8);
  assign w392[42] = |(datain[143:140] ^ 7);
  assign w392[43] = |(datain[139:136] ^ 5);
  assign comp[392] = ~(|w392);
  wire [28-1:0] w393;
  assign w393[0] = |(datain[311:308] ^ 1);
  assign w393[1] = |(datain[307:304] ^ 12);
  assign w393[2] = |(datain[303:300] ^ 2);
  assign w393[3] = |(datain[299:296] ^ 5);
  assign w393[4] = |(datain[295:292] ^ 12);
  assign w393[5] = |(datain[291:288] ^ 13);
  assign w393[6] = |(datain[287:284] ^ 2);
  assign w393[7] = |(datain[283:280] ^ 1);
  assign w393[8] = |(datain[279:276] ^ 11);
  assign w393[9] = |(datain[275:272] ^ 8);
  assign w393[10] = |(datain[271:268] ^ 2);
  assign w393[11] = |(datain[267:264] ^ 1);
  assign w393[12] = |(datain[263:260] ^ 3);
  assign w393[13] = |(datain[259:256] ^ 5);
  assign w393[14] = |(datain[255:252] ^ 12);
  assign w393[15] = |(datain[251:248] ^ 13);
  assign w393[16] = |(datain[247:244] ^ 2);
  assign w393[17] = |(datain[243:240] ^ 1);
  assign w393[18] = |(datain[239:236] ^ 8);
  assign w393[19] = |(datain[235:232] ^ 11);
  assign w393[20] = |(datain[231:228] ^ 13);
  assign w393[21] = |(datain[227:224] ^ 3);
  assign w393[22] = |(datain[223:220] ^ 8);
  assign w393[23] = |(datain[219:216] ^ 13);
  assign w393[24] = |(datain[215:212] ^ 1);
  assign w393[25] = |(datain[211:208] ^ 14);
  assign w393[26] = |(datain[207:204] ^ 2);
  assign w393[27] = |(datain[203:200] ^ 15);
  assign comp[393] = ~(|w393);
  wire [30-1:0] w394;
  assign w394[0] = |(datain[311:308] ^ 9);
  assign w394[1] = |(datain[307:304] ^ 12);
  assign w394[2] = |(datain[303:300] ^ 5);
  assign w394[3] = |(datain[299:296] ^ 0);
  assign w394[4] = |(datain[295:292] ^ 2);
  assign w394[5] = |(datain[291:288] ^ 14);
  assign w394[6] = |(datain[287:284] ^ 10);
  assign w394[7] = |(datain[283:280] ^ 1);
  assign w394[8] = |(datain[279:276] ^ 0);
  assign w394[9] = |(datain[275:272] ^ 7);
  assign w394[10] = |(datain[271:268] ^ 0);
  assign w394[11] = |(datain[267:264] ^ 1);
  assign w394[12] = |(datain[263:260] ^ 4);
  assign w394[13] = |(datain[259:256] ^ 0);
  assign w394[14] = |(datain[255:252] ^ 2);
  assign w394[15] = |(datain[251:248] ^ 14);
  assign w394[16] = |(datain[247:244] ^ 10);
  assign w394[17] = |(datain[243:240] ^ 3);
  assign w394[18] = |(datain[239:236] ^ 0);
  assign w394[19] = |(datain[235:232] ^ 7);
  assign w394[20] = |(datain[231:228] ^ 0);
  assign w394[21] = |(datain[227:224] ^ 1);
  assign w394[22] = |(datain[223:220] ^ 3);
  assign w394[23] = |(datain[219:216] ^ 13);
  assign w394[24] = |(datain[215:212] ^ 0);
  assign w394[25] = |(datain[211:208] ^ 0);
  assign w394[26] = |(datain[207:204] ^ 1);
  assign w394[27] = |(datain[203:200] ^ 0);
  assign w394[28] = |(datain[199:196] ^ 7);
  assign w394[29] = |(datain[195:192] ^ 2);
  assign comp[394] = ~(|w394);
  wire [28-1:0] w395;
  assign w395[0] = |(datain[311:308] ^ 12);
  assign w395[1] = |(datain[307:304] ^ 13);
  assign w395[2] = |(datain[303:300] ^ 7);
  assign w395[3] = |(datain[299:296] ^ 5);
  assign w395[4] = |(datain[295:292] ^ 0);
  assign w395[5] = |(datain[291:288] ^ 3);
  assign w395[6] = |(datain[287:284] ^ 14);
  assign w395[7] = |(datain[283:280] ^ 9);
  assign w395[8] = |(datain[279:276] ^ 12);
  assign w395[9] = |(datain[275:272] ^ 9);
  assign w395[10] = |(datain[271:268] ^ 0);
  assign w395[11] = |(datain[267:264] ^ 0);
  assign w395[12] = |(datain[263:260] ^ 11);
  assign w395[13] = |(datain[259:256] ^ 14);
  assign w395[14] = |(datain[255:252] ^ 0);
  assign w395[15] = |(datain[251:248] ^ 2);
  assign w395[16] = |(datain[247:244] ^ 0);
  assign w395[17] = |(datain[243:240] ^ 0);
  assign w395[18] = |(datain[239:236] ^ 8);
  assign w395[19] = |(datain[235:232] ^ 11);
  assign w395[20] = |(datain[231:228] ^ 0);
  assign w395[21] = |(datain[227:224] ^ 4);
  assign w395[22] = |(datain[223:220] ^ 2);
  assign w395[23] = |(datain[219:216] ^ 13);
  assign w395[24] = |(datain[215:212] ^ 12);
  assign w395[25] = |(datain[211:208] ^ 0);
  assign w395[26] = |(datain[207:204] ^ 0);
  assign w395[27] = |(datain[203:200] ^ 0);
  assign comp[395] = ~(|w395);
  wire [44-1:0] w396;
  assign w396[0] = |(datain[311:308] ^ 2);
  assign w396[1] = |(datain[307:304] ^ 5);
  assign w396[2] = |(datain[303:300] ^ 12);
  assign w396[3] = |(datain[299:296] ^ 13);
  assign w396[4] = |(datain[295:292] ^ 2);
  assign w396[5] = |(datain[291:288] ^ 1);
  assign w396[6] = |(datain[287:284] ^ 0);
  assign w396[7] = |(datain[283:280] ^ 14);
  assign w396[8] = |(datain[279:276] ^ 1);
  assign w396[9] = |(datain[275:272] ^ 15);
  assign w396[10] = |(datain[271:268] ^ 0);
  assign w396[11] = |(datain[267:264] ^ 14);
  assign w396[12] = |(datain[263:260] ^ 0);
  assign w396[13] = |(datain[259:256] ^ 7);
  assign w396[14] = |(datain[255:252] ^ 11);
  assign w396[15] = |(datain[251:248] ^ 4);
  assign w396[16] = |(datain[247:244] ^ 1);
  assign w396[17] = |(datain[243:240] ^ 7);
  assign w396[18] = |(datain[239:236] ^ 9);
  assign w396[19] = |(datain[235:232] ^ 1);
  assign w396[20] = |(datain[231:228] ^ 11);
  assign w396[21] = |(datain[227:224] ^ 4);
  assign w396[22] = |(datain[223:220] ^ 5);
  assign w396[23] = |(datain[219:216] ^ 7);
  assign w396[24] = |(datain[215:212] ^ 2);
  assign w396[25] = |(datain[211:208] ^ 10);
  assign w396[26] = |(datain[207:204] ^ 14);
  assign w396[27] = |(datain[203:200] ^ 5);
  assign w396[28] = |(datain[199:196] ^ 5);
  assign w396[29] = |(datain[195:192] ^ 10);
  assign w396[30] = |(datain[191:188] ^ 5);
  assign w396[31] = |(datain[187:184] ^ 9);
  assign w396[32] = |(datain[183:180] ^ 5);
  assign w396[33] = |(datain[179:176] ^ 11);
  assign w396[34] = |(datain[175:172] ^ 12);
  assign w396[35] = |(datain[171:168] ^ 13);
  assign w396[36] = |(datain[167:164] ^ 0);
  assign w396[37] = |(datain[163:160] ^ 0);
  assign w396[38] = |(datain[159:156] ^ 11);
  assign w396[39] = |(datain[155:152] ^ 4);
  assign w396[40] = |(datain[151:148] ^ 3);
  assign w396[41] = |(datain[147:144] ^ 15);
  assign w396[42] = |(datain[143:140] ^ 11);
  assign w396[43] = |(datain[139:136] ^ 14);
  assign comp[396] = ~(|w396);
  wire [28-1:0] w397;
  assign w397[0] = |(datain[311:308] ^ 2);
  assign w397[1] = |(datain[307:304] ^ 1);
  assign w397[2] = |(datain[303:300] ^ 7);
  assign w397[3] = |(datain[299:296] ^ 2);
  assign w397[4] = |(datain[295:292] ^ 6);
  assign w397[5] = |(datain[291:288] ^ 0);
  assign w397[6] = |(datain[287:284] ^ 11);
  assign w397[7] = |(datain[283:280] ^ 10);
  assign w397[8] = |(datain[279:276] ^ 7);
  assign w397[9] = |(datain[275:272] ^ 13);
  assign w397[10] = |(datain[271:268] ^ 0);
  assign w397[11] = |(datain[267:264] ^ 2);
  assign w397[12] = |(datain[263:260] ^ 11);
  assign w397[13] = |(datain[259:256] ^ 8);
  assign w397[14] = |(datain[255:252] ^ 0);
  assign w397[15] = |(datain[251:248] ^ 2);
  assign w397[16] = |(datain[247:244] ^ 3);
  assign w397[17] = |(datain[243:240] ^ 13);
  assign w397[18] = |(datain[239:236] ^ 12);
  assign w397[19] = |(datain[235:232] ^ 13);
  assign w397[20] = |(datain[231:228] ^ 2);
  assign w397[21] = |(datain[227:224] ^ 1);
  assign w397[22] = |(datain[223:220] ^ 10);
  assign w397[23] = |(datain[219:216] ^ 3);
  assign w397[24] = |(datain[215:212] ^ 1);
  assign w397[25] = |(datain[211:208] ^ 4);
  assign w397[26] = |(datain[207:204] ^ 0);
  assign w397[27] = |(datain[203:200] ^ 1);
  assign comp[397] = ~(|w397);
  wire [28-1:0] w398;
  assign w398[0] = |(datain[311:308] ^ 0);
  assign w398[1] = |(datain[307:304] ^ 14);
  assign w398[2] = |(datain[303:300] ^ 0);
  assign w398[3] = |(datain[299:296] ^ 1);
  assign w398[4] = |(datain[295:292] ^ 0);
  assign w398[5] = |(datain[291:288] ^ 0);
  assign w398[6] = |(datain[287:284] ^ 0);
  assign w398[7] = |(datain[283:280] ^ 0);
  assign w398[8] = |(datain[279:276] ^ 2);
  assign w398[9] = |(datain[275:272] ^ 14);
  assign w398[10] = |(datain[271:268] ^ 8);
  assign w398[11] = |(datain[267:264] ^ 12);
  assign w398[12] = |(datain[263:260] ^ 0);
  assign w398[13] = |(datain[259:256] ^ 6);
  assign w398[14] = |(datain[255:252] ^ 1);
  assign w398[15] = |(datain[251:248] ^ 0);
  assign w398[16] = |(datain[247:244] ^ 0);
  assign w398[17] = |(datain[243:240] ^ 1);
  assign w398[18] = |(datain[239:236] ^ 2);
  assign w398[19] = |(datain[235:232] ^ 14);
  assign w398[20] = |(datain[231:228] ^ 15);
  assign w398[21] = |(datain[227:224] ^ 15);
  assign w398[22] = |(datain[223:220] ^ 2);
  assign w398[23] = |(datain[219:216] ^ 14);
  assign w398[24] = |(datain[215:212] ^ 0);
  assign w398[25] = |(datain[211:208] ^ 14);
  assign w398[26] = |(datain[207:204] ^ 0);
  assign w398[27] = |(datain[203:200] ^ 1);
  assign comp[398] = ~(|w398);
  wire [30-1:0] w399;
  assign w399[0] = |(datain[311:308] ^ 7);
  assign w399[1] = |(datain[307:304] ^ 2);
  assign w399[2] = |(datain[303:300] ^ 5);
  assign w399[3] = |(datain[299:296] ^ 7);
  assign w399[4] = |(datain[295:292] ^ 11);
  assign w399[5] = |(datain[291:288] ^ 10);
  assign w399[6] = |(datain[287:284] ^ 1);
  assign w399[7] = |(datain[283:280] ^ 2);
  assign w399[8] = |(datain[279:276] ^ 0);
  assign w399[9] = |(datain[275:272] ^ 2);
  assign w399[10] = |(datain[271:268] ^ 11);
  assign w399[11] = |(datain[267:264] ^ 8);
  assign w399[12] = |(datain[263:260] ^ 0);
  assign w399[13] = |(datain[259:256] ^ 2);
  assign w399[14] = |(datain[255:252] ^ 3);
  assign w399[15] = |(datain[251:248] ^ 13);
  assign w399[16] = |(datain[247:244] ^ 12);
  assign w399[17] = |(datain[243:240] ^ 13);
  assign w399[18] = |(datain[239:236] ^ 2);
  assign w399[19] = |(datain[235:232] ^ 1);
  assign w399[20] = |(datain[231:228] ^ 10);
  assign w399[21] = |(datain[227:224] ^ 3);
  assign w399[22] = |(datain[223:220] ^ 1);
  assign w399[23] = |(datain[219:216] ^ 4);
  assign w399[24] = |(datain[215:212] ^ 0);
  assign w399[25] = |(datain[211:208] ^ 1);
  assign w399[26] = |(datain[207:204] ^ 8);
  assign w399[27] = |(datain[203:200] ^ 11);
  assign w399[28] = |(datain[199:196] ^ 13);
  assign w399[29] = |(datain[195:192] ^ 8);
  assign comp[399] = ~(|w399);
  wire [46-1:0] w400;
  assign w400[0] = |(datain[311:308] ^ 3);
  assign w400[1] = |(datain[307:304] ^ 15);
  assign w400[2] = |(datain[303:300] ^ 4);
  assign w400[3] = |(datain[299:296] ^ 13);
  assign w400[4] = |(datain[295:292] ^ 5);
  assign w400[5] = |(datain[291:288] ^ 10);
  assign w400[6] = |(datain[287:284] ^ 7);
  assign w400[7] = |(datain[283:280] ^ 4);
  assign w400[8] = |(datain[279:276] ^ 0);
  assign w400[9] = |(datain[275:272] ^ 3);
  assign w400[10] = |(datain[271:268] ^ 14);
  assign w400[11] = |(datain[267:264] ^ 9);
  assign w400[12] = |(datain[263:260] ^ 5);
  assign w400[13] = |(datain[259:256] ^ 3);
  assign w400[14] = |(datain[255:252] ^ 0);
  assign w400[15] = |(datain[251:248] ^ 1);
  assign w400[16] = |(datain[247:244] ^ 14);
  assign w400[17] = |(datain[243:240] ^ 8);
  assign w400[18] = |(datain[239:236] ^ 12);
  assign w400[19] = |(datain[235:232] ^ 9);
  assign w400[20] = |(datain[231:228] ^ 15);
  assign w400[21] = |(datain[227:224] ^ 12);
  assign w400[22] = |(datain[223:220] ^ 12);
  assign w400[23] = |(datain[219:216] ^ 4);
  assign w400[24] = |(datain[215:212] ^ 1);
  assign w400[25] = |(datain[211:208] ^ 14);
  assign w400[26] = |(datain[207:204] ^ 4);
  assign w400[27] = |(datain[203:200] ^ 8);
  assign w400[28] = |(datain[199:196] ^ 0);
  assign w400[29] = |(datain[195:192] ^ 0);
  assign w400[30] = |(datain[191:188] ^ 2);
  assign w400[31] = |(datain[187:184] ^ 6);
  assign w400[32] = |(datain[183:180] ^ 8);
  assign w400[33] = |(datain[179:176] ^ 11);
  assign w400[34] = |(datain[175:172] ^ 4);
  assign w400[35] = |(datain[171:168] ^ 7);
  assign w400[36] = |(datain[167:164] ^ 0);
  assign w400[37] = |(datain[163:160] ^ 15);
  assign w400[38] = |(datain[159:156] ^ 11);
  assign w400[39] = |(datain[155:152] ^ 1);
  assign w400[40] = |(datain[151:148] ^ 0);
  assign w400[41] = |(datain[147:144] ^ 12);
  assign w400[42] = |(datain[143:140] ^ 13);
  assign w400[43] = |(datain[139:136] ^ 3);
  assign w400[44] = |(datain[135:132] ^ 14);
  assign w400[45] = |(datain[131:128] ^ 0);
  assign comp[400] = ~(|w400);
  wire [46-1:0] w401;
  assign w401[0] = |(datain[311:308] ^ 3);
  assign w401[1] = |(datain[307:304] ^ 15);
  assign w401[2] = |(datain[303:300] ^ 4);
  assign w401[3] = |(datain[299:296] ^ 13);
  assign w401[4] = |(datain[295:292] ^ 5);
  assign w401[5] = |(datain[291:288] ^ 10);
  assign w401[6] = |(datain[287:284] ^ 7);
  assign w401[7] = |(datain[283:280] ^ 4);
  assign w401[8] = |(datain[279:276] ^ 0);
  assign w401[9] = |(datain[275:272] ^ 12);
  assign w401[10] = |(datain[271:268] ^ 14);
  assign w401[11] = |(datain[267:264] ^ 8);
  assign w401[12] = |(datain[263:260] ^ 0);
  assign w401[13] = |(datain[259:256] ^ 1);
  assign w401[14] = |(datain[255:252] ^ 0);
  assign w401[15] = |(datain[251:248] ^ 3);
  assign w401[16] = |(datain[247:244] ^ 2);
  assign w401[17] = |(datain[243:240] ^ 11);
  assign w401[18] = |(datain[239:236] ^ 12);
  assign w401[19] = |(datain[235:232] ^ 0);
  assign w401[20] = |(datain[231:228] ^ 5);
  assign w401[21] = |(datain[227:224] ^ 14);
  assign w401[22] = |(datain[223:220] ^ 5);
  assign w401[23] = |(datain[219:216] ^ 15);
  assign w401[24] = |(datain[215:212] ^ 8);
  assign w401[25] = |(datain[211:208] ^ 11);
  assign w401[26] = |(datain[207:204] ^ 14);
  assign w401[27] = |(datain[203:200] ^ 5);
  assign w401[28] = |(datain[199:196] ^ 5);
  assign w401[29] = |(datain[195:192] ^ 13);
  assign w401[30] = |(datain[191:188] ^ 12);
  assign w401[31] = |(datain[187:184] ^ 3);
  assign w401[32] = |(datain[183:180] ^ 9);
  assign w401[33] = |(datain[179:176] ^ 0);
  assign w401[34] = |(datain[175:172] ^ 14);
  assign w401[35] = |(datain[171:168] ^ 8);
  assign w401[36] = |(datain[167:164] ^ 2);
  assign w401[37] = |(datain[163:160] ^ 7);
  assign w401[38] = |(datain[159:156] ^ 0);
  assign w401[39] = |(datain[155:152] ^ 3);
  assign w401[40] = |(datain[151:148] ^ 11);
  assign w401[41] = |(datain[147:144] ^ 1);
  assign w401[42] = |(datain[143:140] ^ 0);
  assign w401[43] = |(datain[139:136] ^ 4);
  assign w401[44] = |(datain[135:132] ^ 12);
  assign w401[45] = |(datain[131:128] ^ 4);
  assign comp[401] = ~(|w401);
  wire [46-1:0] w402;
  assign w402[0] = |(datain[311:308] ^ 11);
  assign w402[1] = |(datain[307:304] ^ 9);
  assign w402[2] = |(datain[303:300] ^ 0);
  assign w402[3] = |(datain[299:296] ^ 1);
  assign w402[4] = |(datain[295:292] ^ 0);
  assign w402[5] = |(datain[291:288] ^ 0);
  assign w402[6] = |(datain[287:284] ^ 13);
  assign w402[7] = |(datain[283:280] ^ 1);
  assign w402[8] = |(datain[279:276] ^ 12);
  assign w402[9] = |(datain[275:272] ^ 2);
  assign w402[10] = |(datain[271:268] ^ 5);
  assign w402[11] = |(datain[267:264] ^ 0);
  assign w402[12] = |(datain[263:260] ^ 12);
  assign w402[13] = |(datain[259:256] ^ 13);
  assign w402[14] = |(datain[255:252] ^ 2);
  assign w402[15] = |(datain[251:248] ^ 6);
  assign w402[16] = |(datain[247:244] ^ 8);
  assign w402[17] = |(datain[243:240] ^ 3);
  assign w402[18] = |(datain[239:236] ^ 12);
  assign w402[19] = |(datain[235:232] ^ 4);
  assign w402[20] = |(datain[231:228] ^ 0);
  assign w402[21] = |(datain[227:224] ^ 2);
  assign w402[22] = |(datain[223:220] ^ 5);
  assign w402[23] = |(datain[219:216] ^ 8);
  assign w402[24] = |(datain[215:212] ^ 5);
  assign w402[25] = |(datain[211:208] ^ 9);
  assign w402[26] = |(datain[207:204] ^ 14);
  assign w402[27] = |(datain[203:200] ^ 2);
  assign w402[28] = |(datain[199:196] ^ 15);
  assign w402[29] = |(datain[195:192] ^ 0);
  assign w402[30] = |(datain[191:188] ^ 15);
  assign w402[31] = |(datain[187:184] ^ 7);
  assign w402[32] = |(datain[183:180] ^ 0);
  assign w402[33] = |(datain[179:176] ^ 6);
  assign w402[34] = |(datain[175:172] ^ 4);
  assign w402[35] = |(datain[171:168] ^ 1);
  assign w402[36] = |(datain[167:164] ^ 0);
  assign w402[37] = |(datain[163:160] ^ 3);
  assign w402[38] = |(datain[159:156] ^ 3);
  assign w402[39] = |(datain[155:152] ^ 15);
  assign w402[40] = |(datain[151:148] ^ 0);
  assign w402[41] = |(datain[147:144] ^ 0);
  assign w402[42] = |(datain[143:140] ^ 7);
  assign w402[43] = |(datain[139:136] ^ 5);
  assign w402[44] = |(datain[135:132] ^ 1);
  assign w402[45] = |(datain[131:128] ^ 1);
  assign comp[402] = ~(|w402);
  wire [48-1:0] w403;
  assign w403[0] = |(datain[311:308] ^ 13);
  assign w403[1] = |(datain[307:304] ^ 12);
  assign w403[2] = |(datain[303:300] ^ 7);
  assign w403[3] = |(datain[299:296] ^ 13);
  assign w403[4] = |(datain[295:292] ^ 4);
  assign w403[5] = |(datain[291:288] ^ 0);
  assign w403[6] = |(datain[287:284] ^ 0);
  assign w403[7] = |(datain[283:280] ^ 2);
  assign w403[8] = |(datain[279:276] ^ 3);
  assign w403[9] = |(datain[275:272] ^ 5);
  assign w403[10] = |(datain[271:268] ^ 5);
  assign w403[11] = |(datain[267:264] ^ 11);
  assign w403[12] = |(datain[263:260] ^ 12);
  assign w403[13] = |(datain[259:256] ^ 3);
  assign w403[14] = |(datain[255:252] ^ 11);
  assign w403[15] = |(datain[251:248] ^ 11);
  assign w403[16] = |(datain[247:244] ^ 11);
  assign w403[17] = |(datain[243:240] ^ 15);
  assign w403[18] = |(datain[239:236] ^ 3);
  assign w403[19] = |(datain[235:232] ^ 5);
  assign w403[20] = |(datain[231:228] ^ 5);
  assign w403[21] = |(datain[227:224] ^ 6);
  assign w403[22] = |(datain[223:220] ^ 6);
  assign w403[23] = |(datain[219:216] ^ 14);
  assign w403[24] = |(datain[215:212] ^ 7);
  assign w403[25] = |(datain[211:208] ^ 8);
  assign w403[26] = |(datain[207:204] ^ 5);
  assign w403[27] = |(datain[203:200] ^ 14);
  assign w403[28] = |(datain[199:196] ^ 2);
  assign w403[29] = |(datain[195:192] ^ 12);
  assign w403[30] = |(datain[191:188] ^ 5);
  assign w403[31] = |(datain[187:184] ^ 9);
  assign w403[32] = |(datain[183:180] ^ 3);
  assign w403[33] = |(datain[179:176] ^ 5);
  assign w403[34] = |(datain[175:172] ^ 4);
  assign w403[35] = |(datain[171:168] ^ 15);
  assign w403[36] = |(datain[167:164] ^ 6);
  assign w403[37] = |(datain[163:160] ^ 3);
  assign w403[38] = |(datain[159:156] ^ 9);
  assign w403[39] = |(datain[155:152] ^ 2);
  assign w403[40] = |(datain[151:148] ^ 3);
  assign w403[41] = |(datain[147:144] ^ 5);
  assign w403[42] = |(datain[143:140] ^ 4);
  assign w403[43] = |(datain[139:136] ^ 11);
  assign w403[44] = |(datain[135:132] ^ 6);
  assign w403[45] = |(datain[131:128] ^ 3);
  assign w403[46] = |(datain[127:124] ^ 8);
  assign w403[47] = |(datain[123:120] ^ 9);
  assign comp[403] = ~(|w403);
  wire [74-1:0] w404;
  assign w404[0] = |(datain[311:308] ^ 2);
  assign w404[1] = |(datain[307:304] ^ 1);
  assign w404[2] = |(datain[303:300] ^ 5);
  assign w404[3] = |(datain[299:296] ^ 9);
  assign w404[4] = |(datain[295:292] ^ 7);
  assign w404[5] = |(datain[291:288] ^ 2);
  assign w404[6] = |(datain[287:284] ^ 2);
  assign w404[7] = |(datain[283:280] ^ 7);
  assign w404[8] = |(datain[279:276] ^ 9);
  assign w404[9] = |(datain[275:272] ^ 7);
  assign w404[10] = |(datain[271:268] ^ 11);
  assign w404[11] = |(datain[267:264] ^ 4);
  assign w404[12] = |(datain[263:260] ^ 4);
  assign w404[13] = |(datain[259:256] ^ 0);
  assign w404[14] = |(datain[255:252] ^ 11);
  assign w404[15] = |(datain[251:248] ^ 11);
  assign w404[16] = |(datain[247:244] ^ 0);
  assign w404[17] = |(datain[243:240] ^ 6);
  assign w404[18] = |(datain[239:236] ^ 0);
  assign w404[19] = |(datain[235:232] ^ 0);
  assign w404[20] = |(datain[231:228] ^ 9);
  assign w404[21] = |(datain[227:224] ^ 9);
  assign w404[22] = |(datain[223:220] ^ 12);
  assign w404[23] = |(datain[219:216] ^ 13);
  assign w404[24] = |(datain[215:212] ^ 2);
  assign w404[25] = |(datain[211:208] ^ 1);
  assign w404[26] = |(datain[207:204] ^ 7);
  assign w404[27] = |(datain[203:200] ^ 2);
  assign w404[28] = |(datain[199:196] ^ 1);
  assign w404[29] = |(datain[195:192] ^ 12);
  assign w404[30] = |(datain[191:188] ^ 3);
  assign w404[31] = |(datain[187:184] ^ 11);
  assign w404[32] = |(datain[183:180] ^ 12);
  assign w404[33] = |(datain[179:176] ^ 1);
  assign w404[34] = |(datain[175:172] ^ 7);
  assign w404[35] = |(datain[171:168] ^ 2);
  assign w404[36] = |(datain[167:164] ^ 1);
  assign w404[37] = |(datain[163:160] ^ 8);
  assign w404[38] = |(datain[159:156] ^ 8);
  assign w404[39] = |(datain[155:152] ^ 3);
  assign w404[40] = |(datain[151:148] ^ 15);
  assign w404[41] = |(datain[147:144] ^ 9);
  assign w404[42] = |(datain[143:140] ^ 15);
  assign w404[43] = |(datain[139:136] ^ 15);
  assign w404[44] = |(datain[135:132] ^ 15);
  assign w404[45] = |(datain[131:128] ^ 8);
  assign w404[46] = |(datain[127:124] ^ 7);
  assign w404[47] = |(datain[123:120] ^ 5);
  assign w404[48] = |(datain[119:116] ^ 1);
  assign w404[49] = |(datain[115:112] ^ 2);
  assign w404[50] = |(datain[111:108] ^ 9);
  assign w404[51] = |(datain[107:104] ^ 7);
  assign w404[52] = |(datain[103:100] ^ 0);
  assign w404[53] = |(datain[99:96] ^ 11);
  assign w404[54] = |(datain[95:92] ^ 12);
  assign w404[55] = |(datain[91:88] ^ 0);
  assign w404[56] = |(datain[87:84] ^ 7);
  assign w404[57] = |(datain[83:80] ^ 4);
  assign w404[58] = |(datain[79:76] ^ 0);
  assign w404[59] = |(datain[75:72] ^ 13);
  assign w404[60] = |(datain[71:68] ^ 11);
  assign w404[61] = |(datain[67:64] ^ 4);
  assign w404[62] = |(datain[63:60] ^ 4);
  assign w404[63] = |(datain[59:56] ^ 0);
  assign w404[64] = |(datain[55:52] ^ 15);
  assign w404[65] = |(datain[51:48] ^ 7);
  assign w404[66] = |(datain[47:44] ^ 13);
  assign w404[67] = |(datain[43:40] ^ 9);
  assign w404[68] = |(datain[39:36] ^ 4);
  assign w404[69] = |(datain[35:32] ^ 10);
  assign w404[70] = |(datain[31:28] ^ 12);
  assign w404[71] = |(datain[27:24] ^ 13);
  assign w404[72] = |(datain[23:20] ^ 2);
  assign w404[73] = |(datain[19:16] ^ 1);
  assign comp[404] = ~(|w404);
  wire [74-1:0] w405;
  assign w405[0] = |(datain[311:308] ^ 5);
  assign w405[1] = |(datain[307:304] ^ 14);
  assign w405[2] = |(datain[303:300] ^ 5);
  assign w405[3] = |(datain[299:296] ^ 11);
  assign w405[4] = |(datain[295:292] ^ 5);
  assign w405[5] = |(datain[291:288] ^ 8);
  assign w405[6] = |(datain[287:284] ^ 0);
  assign w405[7] = |(datain[283:280] ^ 7);
  assign w405[8] = |(datain[279:276] ^ 12);
  assign w405[9] = |(datain[275:272] ^ 3);
  assign w405[10] = |(datain[271:268] ^ 11);
  assign w405[11] = |(datain[267:264] ^ 4);
  assign w405[12] = |(datain[263:260] ^ 3);
  assign w405[13] = |(datain[259:256] ^ 14);
  assign w405[14] = |(datain[255:252] ^ 14);
  assign w405[15] = |(datain[251:248] ^ 11);
  assign w405[16] = |(datain[247:244] ^ 0);
  assign w405[17] = |(datain[243:240] ^ 2);
  assign w405[18] = |(datain[239:236] ^ 11);
  assign w405[19] = |(datain[235:232] ^ 4);
  assign w405[20] = |(datain[231:228] ^ 3);
  assign w405[21] = |(datain[227:224] ^ 15);
  assign w405[22] = |(datain[223:220] ^ 9);
  assign w405[23] = |(datain[219:216] ^ 12);
  assign w405[24] = |(datain[215:212] ^ 2);
  assign w405[25] = |(datain[211:208] ^ 14);
  assign w405[26] = |(datain[207:204] ^ 15);
  assign w405[27] = |(datain[203:200] ^ 15);
  assign w405[28] = |(datain[199:196] ^ 1);
  assign w405[29] = |(datain[195:192] ^ 14);
  assign w405[30] = |(datain[191:188] ^ 15);
  assign w405[31] = |(datain[187:184] ^ 13);
  assign w405[32] = |(datain[183:180] ^ 0);
  assign w405[33] = |(datain[179:176] ^ 4);
  assign w405[34] = |(datain[175:172] ^ 12);
  assign w405[35] = |(datain[171:168] ^ 3);
  assign w405[36] = |(datain[167:164] ^ 3);
  assign w405[37] = |(datain[163:160] ^ 13);
  assign w405[38] = |(datain[159:156] ^ 12);
  assign w405[39] = |(datain[155:152] ^ 13);
  assign w405[40] = |(datain[151:148] ^ 10);
  assign w405[41] = |(datain[147:144] ^ 11);
  assign w405[42] = |(datain[143:140] ^ 7);
  assign w405[43] = |(datain[139:136] ^ 5);
  assign w405[44] = |(datain[135:132] ^ 0);
  assign w405[45] = |(datain[131:128] ^ 7);
  assign w405[46] = |(datain[127:124] ^ 11);
  assign w405[47] = |(datain[123:120] ^ 8);
  assign w405[48] = |(datain[119:116] ^ 15);
  assign w405[49] = |(datain[115:112] ^ 15);
  assign w405[50] = |(datain[111:108] ^ 15);
  assign w405[51] = |(datain[107:104] ^ 15);
  assign w405[52] = |(datain[103:100] ^ 15);
  assign w405[53] = |(datain[99:96] ^ 8);
  assign w405[54] = |(datain[95:92] ^ 12);
  assign w405[55] = |(datain[91:88] ^ 10);
  assign w405[56] = |(datain[87:84] ^ 0);
  assign w405[57] = |(datain[83:80] ^ 2);
  assign w405[58] = |(datain[79:76] ^ 0);
  assign w405[59] = |(datain[75:72] ^ 0);
  assign w405[60] = |(datain[71:68] ^ 3);
  assign w405[61] = |(datain[67:64] ^ 13);
  assign w405[62] = |(datain[63:60] ^ 12);
  assign w405[63] = |(datain[59:56] ^ 0);
  assign w405[64] = |(datain[55:52] ^ 0);
  assign w405[65] = |(datain[51:48] ^ 12);
  assign w405[66] = |(datain[47:44] ^ 7);
  assign w405[67] = |(datain[43:40] ^ 5);
  assign w405[68] = |(datain[39:36] ^ 0);
  assign w405[69] = |(datain[35:32] ^ 3);
  assign w405[70] = |(datain[31:28] ^ 8);
  assign w405[71] = |(datain[27:24] ^ 6);
  assign w405[72] = |(datain[23:20] ^ 12);
  assign w405[73] = |(datain[19:16] ^ 4);
  assign comp[405] = ~(|w405);
  wire [30-1:0] w406;
  assign w406[0] = |(datain[311:308] ^ 1);
  assign w406[1] = |(datain[307:304] ^ 9);
  assign w406[2] = |(datain[303:300] ^ 0);
  assign w406[3] = |(datain[299:296] ^ 0);
  assign w406[4] = |(datain[295:292] ^ 0);
  assign w406[5] = |(datain[291:288] ^ 14);
  assign w406[6] = |(datain[287:284] ^ 1);
  assign w406[7] = |(datain[283:280] ^ 15);
  assign w406[8] = |(datain[279:276] ^ 11);
  assign w406[9] = |(datain[275:272] ^ 10);
  assign w406[10] = |(datain[271:268] ^ 5);
  assign w406[11] = |(datain[267:264] ^ 12);
  assign w406[12] = |(datain[263:260] ^ 0);
  assign w406[13] = |(datain[259:256] ^ 2);
  assign w406[14] = |(datain[255:252] ^ 11);
  assign w406[15] = |(datain[251:248] ^ 8);
  assign w406[16] = |(datain[247:244] ^ 2);
  assign w406[17] = |(datain[243:240] ^ 1);
  assign w406[18] = |(datain[239:236] ^ 2);
  assign w406[19] = |(datain[235:232] ^ 5);
  assign w406[20] = |(datain[231:228] ^ 12);
  assign w406[21] = |(datain[227:224] ^ 13);
  assign w406[22] = |(datain[223:220] ^ 2);
  assign w406[23] = |(datain[219:216] ^ 1);
  assign w406[24] = |(datain[215:212] ^ 8);
  assign w406[25] = |(datain[211:208] ^ 14);
  assign w406[26] = |(datain[207:204] ^ 0);
  assign w406[27] = |(datain[203:200] ^ 6);
  assign w406[28] = |(datain[199:196] ^ 3);
  assign w406[29] = |(datain[195:192] ^ 1);
  assign comp[406] = ~(|w406);
  wire [44-1:0] w407;
  assign w407[0] = |(datain[311:308] ^ 12);
  assign w407[1] = |(datain[307:304] ^ 13);
  assign w407[2] = |(datain[303:300] ^ 2);
  assign w407[3] = |(datain[299:296] ^ 1);
  assign w407[4] = |(datain[295:292] ^ 8);
  assign w407[5] = |(datain[291:288] ^ 0);
  assign w407[6] = |(datain[287:284] ^ 15);
  assign w407[7] = |(datain[283:280] ^ 12);
  assign w407[8] = |(datain[279:276] ^ 14);
  assign w407[9] = |(datain[275:272] ^ 1);
  assign w407[10] = |(datain[271:268] ^ 7);
  assign w407[11] = |(datain[267:264] ^ 3);
  assign w407[12] = |(datain[263:260] ^ 1);
  assign w407[13] = |(datain[259:256] ^ 3);
  assign w407[14] = |(datain[255:252] ^ 8);
  assign w407[15] = |(datain[251:248] ^ 0);
  assign w407[16] = |(datain[247:244] ^ 15);
  assign w407[17] = |(datain[243:240] ^ 12);
  assign w407[18] = |(datain[239:236] ^ 0);
  assign w407[19] = |(datain[235:232] ^ 3);
  assign w407[20] = |(datain[231:228] ^ 0);
  assign w407[21] = |(datain[227:224] ^ 7);
  assign w407[22] = |(datain[223:220] ^ 2);
  assign w407[23] = |(datain[219:216] ^ 14);
  assign w407[24] = |(datain[215:212] ^ 8);
  assign w407[25] = |(datain[211:208] ^ 14);
  assign w407[26] = |(datain[207:204] ^ 1);
  assign w407[27] = |(datain[203:200] ^ 6);
  assign w407[28] = |(datain[199:196] ^ 4);
  assign w407[29] = |(datain[195:192] ^ 5);
  assign w407[30] = |(datain[191:188] ^ 0);
  assign w407[31] = |(datain[187:184] ^ 0);
  assign w407[32] = |(datain[183:180] ^ 2);
  assign w407[33] = |(datain[179:176] ^ 14);
  assign w407[34] = |(datain[175:172] ^ 8);
  assign w407[35] = |(datain[171:168] ^ 11);
  assign w407[36] = |(datain[167:164] ^ 2);
  assign w407[37] = |(datain[163:160] ^ 6);
  assign w407[38] = |(datain[159:156] ^ 4);
  assign w407[39] = |(datain[155:152] ^ 3);
  assign w407[40] = |(datain[151:148] ^ 0);
  assign w407[41] = |(datain[147:144] ^ 0);
  assign w407[42] = |(datain[143:140] ^ 2);
  assign w407[43] = |(datain[139:136] ^ 14);
  assign comp[407] = ~(|w407);
  wire [76-1:0] w408;
  assign w408[0] = |(datain[311:308] ^ 2);
  assign w408[1] = |(datain[307:304] ^ 14);
  assign w408[2] = |(datain[303:300] ^ 10);
  assign w408[3] = |(datain[299:296] ^ 3);
  assign w408[4] = |(datain[295:292] ^ 0);
  assign w408[5] = |(datain[291:288] ^ 5);
  assign w408[6] = |(datain[287:284] ^ 0);
  assign w408[7] = |(datain[283:280] ^ 1);
  assign w408[8] = |(datain[279:276] ^ 14);
  assign w408[9] = |(datain[275:272] ^ 8);
  assign w408[10] = |(datain[271:268] ^ 2);
  assign w408[11] = |(datain[267:264] ^ 3);
  assign w408[12] = |(datain[263:260] ^ 0);
  assign w408[13] = |(datain[259:256] ^ 1);
  assign w408[14] = |(datain[255:252] ^ 8);
  assign w408[15] = |(datain[251:248] ^ 13);
  assign w408[16] = |(datain[247:244] ^ 1);
  assign w408[17] = |(datain[243:240] ^ 6);
  assign w408[18] = |(datain[239:236] ^ 0);
  assign w408[19] = |(datain[235:232] ^ 4);
  assign w408[20] = |(datain[231:228] ^ 0);
  assign w408[21] = |(datain[227:224] ^ 1);
  assign w408[22] = |(datain[223:220] ^ 11);
  assign w408[23] = |(datain[219:216] ^ 9);
  assign w408[24] = |(datain[215:212] ^ 0);
  assign w408[25] = |(datain[211:208] ^ 3);
  assign w408[26] = |(datain[207:204] ^ 0);
  assign w408[27] = |(datain[203:200] ^ 0);
  assign w408[28] = |(datain[199:196] ^ 11);
  assign w408[29] = |(datain[195:192] ^ 4);
  assign w408[30] = |(datain[191:188] ^ 4);
  assign w408[31] = |(datain[187:184] ^ 0);
  assign w408[32] = |(datain[183:180] ^ 12);
  assign w408[33] = |(datain[179:176] ^ 13);
  assign w408[34] = |(datain[175:172] ^ 2);
  assign w408[35] = |(datain[171:168] ^ 1);
  assign w408[36] = |(datain[167:164] ^ 7);
  assign w408[37] = |(datain[163:160] ^ 2);
  assign w408[38] = |(datain[159:156] ^ 2);
  assign w408[39] = |(datain[155:152] ^ 10);
  assign w408[40] = |(datain[151:148] ^ 3);
  assign w408[41] = |(datain[147:144] ^ 3);
  assign w408[42] = |(datain[143:140] ^ 13);
  assign w408[43] = |(datain[139:136] ^ 2);
  assign w408[44] = |(datain[135:132] ^ 2);
  assign w408[45] = |(datain[131:128] ^ 14);
  assign w408[46] = |(datain[127:124] ^ 8);
  assign w408[47] = |(datain[123:120] ^ 9);
  assign w408[48] = |(datain[119:116] ^ 1);
  assign w408[49] = |(datain[115:112] ^ 6);
  assign w408[50] = |(datain[111:108] ^ 1);
  assign w408[51] = |(datain[107:104] ^ 12);
  assign w408[52] = |(datain[103:100] ^ 0);
  assign w408[53] = |(datain[99:96] ^ 1);
  assign w408[54] = |(datain[95:92] ^ 14);
  assign w408[55] = |(datain[91:88] ^ 8);
  assign w408[56] = |(datain[87:84] ^ 1);
  assign w408[57] = |(datain[83:80] ^ 6);
  assign w408[58] = |(datain[79:76] ^ 0);
  assign w408[59] = |(datain[75:72] ^ 1);
  assign w408[60] = |(datain[71:68] ^ 14);
  assign w408[61] = |(datain[67:64] ^ 8);
  assign w408[62] = |(datain[63:60] ^ 14);
  assign w408[63] = |(datain[59:56] ^ 2);
  assign w408[64] = |(datain[55:52] ^ 0);
  assign w408[65] = |(datain[51:48] ^ 0);
  assign w408[66] = |(datain[47:44] ^ 2);
  assign w408[67] = |(datain[43:40] ^ 14);
  assign w408[68] = |(datain[39:36] ^ 8);
  assign w408[69] = |(datain[35:32] ^ 11);
  assign w408[70] = |(datain[31:28] ^ 0);
  assign w408[71] = |(datain[27:24] ^ 14);
  assign w408[72] = |(datain[23:20] ^ 6);
  assign w408[73] = |(datain[19:16] ^ 10);
  assign w408[74] = |(datain[15:12] ^ 0);
  assign w408[75] = |(datain[11:8] ^ 5);
  assign comp[408] = ~(|w408);
  wire [74-1:0] w409;
  assign w409[0] = |(datain[311:308] ^ 7);
  assign w409[1] = |(datain[307:304] ^ 6);
  assign w409[2] = |(datain[303:300] ^ 2);
  assign w409[3] = |(datain[299:296] ^ 4);
  assign w409[4] = |(datain[295:292] ^ 11);
  assign w409[5] = |(datain[291:288] ^ 0);
  assign w409[6] = |(datain[287:284] ^ 0);
  assign w409[7] = |(datain[283:280] ^ 2);
  assign w409[8] = |(datain[279:276] ^ 11);
  assign w409[9] = |(datain[275:272] ^ 9);
  assign w409[10] = |(datain[271:268] ^ 0);
  assign w409[11] = |(datain[267:264] ^ 1);
  assign w409[12] = |(datain[263:260] ^ 0);
  assign w409[13] = |(datain[259:256] ^ 0);
  assign w409[14] = |(datain[255:252] ^ 3);
  assign w409[15] = |(datain[251:248] ^ 3);
  assign w409[16] = |(datain[247:244] ^ 13);
  assign w409[17] = |(datain[243:240] ^ 2);
  assign w409[18] = |(datain[239:236] ^ 8);
  assign w409[19] = |(datain[235:232] ^ 1);
  assign w409[20] = |(datain[231:228] ^ 12);
  assign w409[21] = |(datain[227:224] ^ 3);
  assign w409[22] = |(datain[223:220] ^ 5);
  assign w409[23] = |(datain[219:216] ^ 3);
  assign w409[24] = |(datain[215:212] ^ 0);
  assign w409[25] = |(datain[211:208] ^ 3);
  assign w409[26] = |(datain[207:204] ^ 8);
  assign w409[27] = |(datain[203:200] ^ 11);
  assign w409[28] = |(datain[199:196] ^ 15);
  assign w409[29] = |(datain[195:192] ^ 3);
  assign w409[30] = |(datain[191:188] ^ 0);
  assign w409[31] = |(datain[187:184] ^ 14);
  assign w409[32] = |(datain[183:180] ^ 1);
  assign w409[33] = |(datain[179:176] ^ 15);
  assign w409[34] = |(datain[175:172] ^ 12);
  assign w409[35] = |(datain[171:168] ^ 13);
  assign w409[36] = |(datain[167:164] ^ 2);
  assign w409[37] = |(datain[163:160] ^ 5);
  assign w409[38] = |(datain[159:156] ^ 7);
  assign w409[39] = |(datain[155:152] ^ 2);
  assign w409[40] = |(datain[151:148] ^ 1);
  assign w409[41] = |(datain[147:144] ^ 0);
  assign w409[42] = |(datain[143:140] ^ 9);
  assign w409[43] = |(datain[139:136] ^ 13);
  assign w409[44] = |(datain[135:132] ^ 11);
  assign w409[45] = |(datain[131:128] ^ 0);
  assign w409[46] = |(datain[127:124] ^ 0);
  assign w409[47] = |(datain[123:120] ^ 2);
  assign w409[48] = |(datain[119:116] ^ 8);
  assign w409[49] = |(datain[115:112] ^ 11);
  assign w409[50] = |(datain[111:108] ^ 13);
  assign w409[51] = |(datain[107:104] ^ 14);
  assign w409[52] = |(datain[103:100] ^ 11);
  assign w409[53] = |(datain[99:96] ^ 9);
  assign w409[54] = |(datain[95:92] ^ 0);
  assign w409[55] = |(datain[91:88] ^ 1);
  assign w409[56] = |(datain[87:84] ^ 0);
  assign w409[57] = |(datain[83:80] ^ 0);
  assign w409[58] = |(datain[79:76] ^ 3);
  assign w409[59] = |(datain[75:72] ^ 3);
  assign w409[60] = |(datain[71:68] ^ 13);
  assign w409[61] = |(datain[67:64] ^ 2);
  assign w409[62] = |(datain[63:60] ^ 12);
  assign w409[63] = |(datain[59:56] ^ 6);
  assign w409[64] = |(datain[55:52] ^ 4);
  assign w409[65] = |(datain[51:48] ^ 4);
  assign w409[66] = |(datain[47:44] ^ 1);
  assign w409[67] = |(datain[43:40] ^ 10);
  assign w409[68] = |(datain[39:36] ^ 0);
  assign w409[69] = |(datain[35:32] ^ 0);
  assign w409[70] = |(datain[31:28] ^ 12);
  assign w409[71] = |(datain[27:24] ^ 13);
  assign w409[72] = |(datain[23:20] ^ 2);
  assign w409[73] = |(datain[19:16] ^ 6);
  assign comp[409] = ~(|w409);
  wire [46-1:0] w410;
  assign w410[0] = |(datain[311:308] ^ 0);
  assign w410[1] = |(datain[307:304] ^ 8);
  assign w410[2] = |(datain[303:300] ^ 0);
  assign w410[3] = |(datain[299:296] ^ 1);
  assign w410[4] = |(datain[295:292] ^ 2);
  assign w410[5] = |(datain[291:288] ^ 6);
  assign w410[6] = |(datain[287:284] ^ 10);
  assign w410[7] = |(datain[283:280] ^ 3);
  assign w410[8] = |(datain[279:276] ^ 8);
  assign w410[9] = |(datain[275:272] ^ 6);
  assign w410[10] = |(datain[271:268] ^ 0);
  assign w410[11] = |(datain[267:264] ^ 0);
  assign w410[12] = |(datain[263:260] ^ 2);
  assign w410[13] = |(datain[259:256] ^ 6);
  assign w410[14] = |(datain[255:252] ^ 12);
  assign w410[15] = |(datain[251:248] ^ 7);
  assign w410[16] = |(datain[247:244] ^ 0);
  assign w410[17] = |(datain[243:240] ^ 6);
  assign w410[18] = |(datain[239:236] ^ 8);
  assign w410[19] = |(datain[235:232] ^ 4);
  assign w410[20] = |(datain[231:228] ^ 0);
  assign w410[21] = |(datain[227:224] ^ 0);
  assign w410[22] = |(datain[223:220] ^ 7);
  assign w410[23] = |(datain[219:216] ^ 3);
  assign w410[24] = |(datain[215:212] ^ 0);
  assign w410[25] = |(datain[211:208] ^ 1);
  assign w410[26] = |(datain[207:204] ^ 2);
  assign w410[27] = |(datain[203:200] ^ 6);
  assign w410[28] = |(datain[199:196] ^ 10);
  assign w410[29] = |(datain[195:192] ^ 3);
  assign w410[30] = |(datain[191:188] ^ 7);
  assign w410[31] = |(datain[187:184] ^ 2);
  assign w410[32] = |(datain[183:180] ^ 0);
  assign w410[33] = |(datain[179:176] ^ 0);
  assign w410[34] = |(datain[175:172] ^ 2);
  assign w410[35] = |(datain[171:168] ^ 6);
  assign w410[36] = |(datain[167:164] ^ 12);
  assign w410[37] = |(datain[163:160] ^ 7);
  assign w410[38] = |(datain[159:156] ^ 0);
  assign w410[39] = |(datain[155:152] ^ 6);
  assign w410[40] = |(datain[151:148] ^ 7);
  assign w410[41] = |(datain[147:144] ^ 0);
  assign w410[42] = |(datain[143:140] ^ 0);
  assign w410[43] = |(datain[139:136] ^ 0);
  assign w410[44] = |(datain[135:132] ^ 11);
  assign w410[45] = |(datain[131:128] ^ 13);
  assign comp[410] = ~(|w410);
  wire [44-1:0] w411;
  assign w411[0] = |(datain[311:308] ^ 5);
  assign w411[1] = |(datain[307:304] ^ 3);
  assign w411[2] = |(datain[303:300] ^ 8);
  assign w411[3] = |(datain[299:296] ^ 0);
  assign w411[4] = |(datain[295:292] ^ 7);
  assign w411[5] = |(datain[291:288] ^ 7);
  assign w411[6] = |(datain[287:284] ^ 1);
  assign w411[7] = |(datain[283:280] ^ 0);
  assign w411[8] = |(datain[279:276] ^ 13);
  assign w411[9] = |(datain[275:272] ^ 14);
  assign w411[10] = |(datain[271:268] ^ 9);
  assign w411[11] = |(datain[267:264] ^ 0);
  assign w411[12] = |(datain[263:260] ^ 11);
  assign w411[13] = |(datain[259:256] ^ 9);
  assign w411[14] = |(datain[255:252] ^ 15);
  assign w411[15] = |(datain[251:248] ^ 2);
  assign w411[16] = |(datain[247:244] ^ 0);
  assign w411[17] = |(datain[243:240] ^ 3);
  assign w411[18] = |(datain[239:236] ^ 8);
  assign w411[19] = |(datain[235:232] ^ 3);
  assign w411[20] = |(datain[231:228] ^ 12);
  assign w411[21] = |(datain[227:224] ^ 3);
  assign w411[22] = |(datain[223:220] ^ 1);
  assign w411[23] = |(datain[219:216] ^ 15);
  assign w411[24] = |(datain[215:212] ^ 9);
  assign w411[25] = |(datain[211:208] ^ 0);
  assign w411[26] = |(datain[207:204] ^ 8);
  assign w411[27] = |(datain[203:200] ^ 10);
  assign w411[28] = |(datain[199:196] ^ 0);
  assign w411[29] = |(datain[195:192] ^ 7);
  assign w411[30] = |(datain[191:188] ^ 3);
  assign w411[31] = |(datain[187:184] ^ 4);
  assign w411[32] = |(datain[183:180] ^ 3);
  assign w411[33] = |(datain[179:176] ^ 10);
  assign w411[34] = |(datain[175:172] ^ 8);
  assign w411[35] = |(datain[171:168] ^ 8);
  assign w411[36] = |(datain[167:164] ^ 0);
  assign w411[37] = |(datain[163:160] ^ 7);
  assign w411[38] = |(datain[159:156] ^ 4);
  assign w411[39] = |(datain[155:152] ^ 3);
  assign w411[40] = |(datain[151:148] ^ 14);
  assign w411[41] = |(datain[147:144] ^ 2);
  assign w411[42] = |(datain[143:140] ^ 15);
  assign w411[43] = |(datain[139:136] ^ 7);
  assign comp[411] = ~(|w411);
  wire [46-1:0] w412;
  assign w412[0] = |(datain[311:308] ^ 8);
  assign w412[1] = |(datain[307:304] ^ 10);
  assign w412[2] = |(datain[303:300] ^ 9);
  assign w412[3] = |(datain[299:296] ^ 14);
  assign w412[4] = |(datain[295:292] ^ 1);
  assign w412[5] = |(datain[291:288] ^ 4);
  assign w412[6] = |(datain[287:284] ^ 0);
  assign w412[7] = |(datain[283:280] ^ 1);
  assign w412[8] = |(datain[279:276] ^ 11);
  assign w412[9] = |(datain[275:272] ^ 15);
  assign w412[10] = |(datain[271:268] ^ 10);
  assign w412[11] = |(datain[267:264] ^ 15);
  assign w412[12] = |(datain[263:260] ^ 0);
  assign w412[13] = |(datain[259:256] ^ 3);
  assign w412[14] = |(datain[255:252] ^ 8);
  assign w412[15] = |(datain[251:248] ^ 11);
  assign w412[16] = |(datain[247:244] ^ 12);
  assign w412[17] = |(datain[243:240] ^ 15);
  assign w412[18] = |(datain[239:236] ^ 8);
  assign w412[19] = |(datain[235:232] ^ 13);
  assign w412[20] = |(datain[231:228] ^ 11);
  assign w412[21] = |(datain[227:224] ^ 6);
  assign w412[22] = |(datain[223:220] ^ 2);
  assign w412[23] = |(datain[219:216] ^ 13);
  assign w412[24] = |(datain[215:212] ^ 0);
  assign w412[25] = |(datain[211:208] ^ 1);
  assign w412[26] = |(datain[207:204] ^ 2);
  assign w412[27] = |(datain[203:200] ^ 14);
  assign w412[28] = |(datain[199:196] ^ 3);
  assign w412[29] = |(datain[195:192] ^ 0);
  assign w412[30] = |(datain[191:188] ^ 1);
  assign w412[31] = |(datain[187:184] ^ 12);
  assign w412[32] = |(datain[183:180] ^ 4);
  assign w412[33] = |(datain[179:176] ^ 6);
  assign w412[34] = |(datain[175:172] ^ 11);
  assign w412[35] = |(datain[171:168] ^ 4);
  assign w412[36] = |(datain[167:164] ^ 2);
  assign w412[37] = |(datain[163:160] ^ 14);
  assign w412[38] = |(datain[159:156] ^ 12);
  assign w412[39] = |(datain[155:152] ^ 13);
  assign w412[40] = |(datain[151:148] ^ 2);
  assign w412[41] = |(datain[147:144] ^ 1);
  assign w412[42] = |(datain[143:140] ^ 14);
  assign w412[43] = |(datain[139:136] ^ 0);
  assign w412[44] = |(datain[135:132] ^ 15);
  assign w412[45] = |(datain[131:128] ^ 6);
  assign comp[412] = ~(|w412);
  wire [42-1:0] w413;
  assign w413[0] = |(datain[311:308] ^ 2);
  assign w413[1] = |(datain[307:304] ^ 14);
  assign w413[2] = |(datain[303:300] ^ 8);
  assign w413[3] = |(datain[299:296] ^ 10);
  assign w413[4] = |(datain[295:292] ^ 0);
  assign w413[5] = |(datain[291:288] ^ 4);
  assign w413[6] = |(datain[287:284] ^ 3);
  assign w413[7] = |(datain[283:280] ^ 2);
  assign w413[8] = |(datain[279:276] ^ 12);
  assign w413[9] = |(datain[275:272] ^ 4);
  assign w413[10] = |(datain[271:268] ^ 2);
  assign w413[11] = |(datain[267:264] ^ 14);
  assign w413[12] = |(datain[263:260] ^ 8);
  assign w413[13] = |(datain[259:256] ^ 8);
  assign w413[14] = |(datain[255:252] ^ 0);
  assign w413[15] = |(datain[251:248] ^ 4);
  assign w413[16] = |(datain[247:244] ^ 4);
  assign w413[17] = |(datain[243:240] ^ 6);
  assign w413[18] = |(datain[239:236] ^ 3);
  assign w413[19] = |(datain[235:232] ^ 11);
  assign w413[20] = |(datain[231:228] ^ 15);
  assign w413[21] = |(datain[227:224] ^ 1);
  assign w413[22] = |(datain[223:220] ^ 7);
  assign w413[23] = |(datain[219:216] ^ 5);
  assign w413[24] = |(datain[215:212] ^ 15);
  assign w413[25] = |(datain[211:208] ^ 3);
  assign w413[26] = |(datain[207:204] ^ 12);
  assign w413[27] = |(datain[203:200] ^ 3);
  assign w413[28] = |(datain[199:196] ^ 11);
  assign w413[29] = |(datain[195:192] ^ 4);
  assign w413[30] = |(datain[191:188] ^ 2);
  assign w413[31] = |(datain[187:184] ^ 12);
  assign w413[32] = |(datain[183:180] ^ 12);
  assign w413[33] = |(datain[179:176] ^ 13);
  assign w413[34] = |(datain[175:172] ^ 2);
  assign w413[35] = |(datain[171:168] ^ 1);
  assign w413[36] = |(datain[167:164] ^ 0);
  assign w413[37] = |(datain[163:160] ^ 2);
  assign w413[38] = |(datain[159:156] ^ 12);
  assign w413[39] = |(datain[155:152] ^ 4);
  assign w413[40] = |(datain[151:148] ^ 0);
  assign w413[41] = |(datain[147:144] ^ 2);
  assign comp[413] = ~(|w413);
  wire [74-1:0] w414;
  assign w414[0] = |(datain[311:308] ^ 2);
  assign w414[1] = |(datain[307:304] ^ 10);
  assign w414[2] = |(datain[303:300] ^ 12);
  assign w414[3] = |(datain[299:296] ^ 13);
  assign w414[4] = |(datain[295:292] ^ 2);
  assign w414[5] = |(datain[291:288] ^ 1);
  assign w414[6] = |(datain[287:284] ^ 3);
  assign w414[7] = |(datain[283:280] ^ 12);
  assign w414[8] = |(datain[279:276] ^ 0);
  assign w414[9] = |(datain[275:272] ^ 1);
  assign w414[10] = |(datain[271:268] ^ 7);
  assign w414[11] = |(datain[267:264] ^ 4);
  assign w414[12] = |(datain[263:260] ^ 0);
  assign w414[13] = |(datain[259:256] ^ 14);
  assign w414[14] = |(datain[255:252] ^ 3);
  assign w414[15] = |(datain[251:248] ^ 12);
  assign w414[16] = |(datain[247:244] ^ 0);
  assign w414[17] = |(datain[243:240] ^ 3);
  assign w414[18] = |(datain[239:236] ^ 7);
  assign w414[19] = |(datain[235:232] ^ 4);
  assign w414[20] = |(datain[231:228] ^ 0);
  assign w414[21] = |(datain[227:224] ^ 10);
  assign w414[22] = |(datain[223:220] ^ 3);
  assign w414[23] = |(datain[219:216] ^ 12);
  assign w414[24] = |(datain[215:212] ^ 0);
  assign w414[25] = |(datain[211:208] ^ 5);
  assign w414[26] = |(datain[207:204] ^ 7);
  assign w414[27] = |(datain[203:200] ^ 4);
  assign w414[28] = |(datain[199:196] ^ 0);
  assign w414[29] = |(datain[195:192] ^ 6);
  assign w414[30] = |(datain[191:188] ^ 14);
  assign w414[31] = |(datain[187:184] ^ 8);
  assign w414[32] = |(datain[183:180] ^ 2);
  assign w414[33] = |(datain[179:176] ^ 4);
  assign w414[34] = |(datain[175:172] ^ 0);
  assign w414[35] = |(datain[171:168] ^ 3);
  assign w414[36] = |(datain[167:164] ^ 14);
  assign w414[37] = |(datain[163:160] ^ 11);
  assign w414[38] = |(datain[159:156] ^ 0);
  assign w414[39] = |(datain[155:152] ^ 4);
  assign w414[40] = |(datain[151:148] ^ 9);
  assign w414[41] = |(datain[147:144] ^ 0);
  assign w414[42] = |(datain[143:140] ^ 14);
  assign w414[43] = |(datain[139:136] ^ 8);
  assign w414[44] = |(datain[135:132] ^ 1);
  assign w414[45] = |(datain[131:128] ^ 7);
  assign w414[46] = |(datain[127:124] ^ 0);
  assign w414[47] = |(datain[123:120] ^ 3);
  assign w414[48] = |(datain[119:116] ^ 11);
  assign w414[49] = |(datain[115:112] ^ 14);
  assign w414[50] = |(datain[111:108] ^ 13);
  assign w414[51] = |(datain[107:104] ^ 15);
  assign w414[52] = |(datain[103:100] ^ 10);
  assign w414[53] = |(datain[99:96] ^ 15);
  assign w414[54] = |(datain[95:92] ^ 11);
  assign w414[55] = |(datain[91:88] ^ 4);
  assign w414[56] = |(datain[87:84] ^ 3);
  assign w414[57] = |(datain[83:80] ^ 0);
  assign w414[58] = |(datain[79:76] ^ 12);
  assign w414[59] = |(datain[75:72] ^ 13);
  assign w414[60] = |(datain[71:68] ^ 2);
  assign w414[61] = |(datain[67:64] ^ 1);
  assign w414[62] = |(datain[63:60] ^ 8);
  assign w414[63] = |(datain[59:56] ^ 1);
  assign w414[64] = |(datain[55:52] ^ 15);
  assign w414[65] = |(datain[51:48] ^ 15);
  assign w414[66] = |(datain[47:44] ^ 12);
  assign w414[67] = |(datain[43:40] ^ 3);
  assign w414[68] = |(datain[39:36] ^ 12);
  assign w414[69] = |(datain[35:32] ^ 3);
  assign w414[70] = |(datain[31:28] ^ 7);
  assign w414[71] = |(datain[27:24] ^ 5);
  assign w414[72] = |(datain[23:20] ^ 1);
  assign w414[73] = |(datain[19:16] ^ 12);
  assign comp[414] = ~(|w414);
  wire [42-1:0] w415;
  assign w415[0] = |(datain[311:308] ^ 0);
  assign w415[1] = |(datain[307:304] ^ 3);
  assign w415[2] = |(datain[303:300] ^ 14);
  assign w415[3] = |(datain[299:296] ^ 9);
  assign w415[4] = |(datain[295:292] ^ 11);
  assign w415[5] = |(datain[291:288] ^ 3);
  assign w415[6] = |(datain[287:284] ^ 15);
  assign w415[7] = |(datain[283:280] ^ 13);
  assign w415[8] = |(datain[279:276] ^ 8);
  assign w415[9] = |(datain[275:272] ^ 0);
  assign w415[10] = |(datain[271:268] ^ 15);
  assign w415[11] = |(datain[267:264] ^ 12);
  assign w415[12] = |(datain[263:260] ^ 3);
  assign w415[13] = |(datain[259:256] ^ 0);
  assign w415[14] = |(datain[255:252] ^ 7);
  assign w415[15] = |(datain[251:248] ^ 5);
  assign w415[16] = |(datain[247:244] ^ 0);
  assign w415[17] = |(datain[243:240] ^ 9);
  assign w415[18] = |(datain[239:236] ^ 8);
  assign w415[19] = |(datain[235:232] ^ 1);
  assign w415[20] = |(datain[231:228] ^ 15);
  assign w415[21] = |(datain[227:224] ^ 14);
  assign w415[22] = |(datain[223:220] ^ 10);
  assign w415[23] = |(datain[219:216] ^ 3);
  assign w415[24] = |(datain[215:212] ^ 11);
  assign w415[25] = |(datain[211:208] ^ 4);
  assign w415[26] = |(datain[207:204] ^ 7);
  assign w415[27] = |(datain[203:200] ^ 5);
  assign w415[28] = |(datain[199:196] ^ 0);
  assign w415[29] = |(datain[195:192] ^ 3);
  assign w415[30] = |(datain[191:188] ^ 11);
  assign w415[31] = |(datain[187:184] ^ 15);
  assign w415[32] = |(datain[183:180] ^ 12);
  assign w415[33] = |(datain[179:176] ^ 10);
  assign w415[34] = |(datain[175:172] ^ 11);
  assign w415[35] = |(datain[171:168] ^ 13);
  assign w415[36] = |(datain[167:164] ^ 15);
  assign w415[37] = |(datain[163:160] ^ 11);
  assign w415[38] = |(datain[159:156] ^ 2);
  assign w415[39] = |(datain[155:152] ^ 14);
  assign w415[40] = |(datain[151:148] ^ 15);
  assign w415[41] = |(datain[147:144] ^ 15);
  assign comp[415] = ~(|w415);
  wire [44-1:0] w416;
  assign w416[0] = |(datain[311:308] ^ 15);
  assign w416[1] = |(datain[307:304] ^ 12);
  assign w416[2] = |(datain[303:300] ^ 4);
  assign w416[3] = |(datain[299:296] ^ 11);
  assign w416[4] = |(datain[295:292] ^ 7);
  assign w416[5] = |(datain[291:288] ^ 5);
  assign w416[6] = |(datain[287:284] ^ 0);
  assign w416[7] = |(datain[283:280] ^ 3);
  assign w416[8] = |(datain[279:276] ^ 14);
  assign w416[9] = |(datain[275:272] ^ 9);
  assign w416[10] = |(datain[271:268] ^ 8);
  assign w416[11] = |(datain[267:264] ^ 13);
  assign w416[12] = |(datain[263:260] ^ 15);
  assign w416[13] = |(datain[259:256] ^ 13);
  assign w416[14] = |(datain[255:252] ^ 8);
  assign w416[15] = |(datain[251:248] ^ 0);
  assign w416[16] = |(datain[247:244] ^ 15);
  assign w416[17] = |(datain[243:240] ^ 12);
  assign w416[18] = |(datain[239:236] ^ 3);
  assign w416[19] = |(datain[235:232] ^ 0);
  assign w416[20] = |(datain[231:228] ^ 7);
  assign w416[21] = |(datain[227:224] ^ 5);
  assign w416[22] = |(datain[223:220] ^ 0);
  assign w416[23] = |(datain[219:216] ^ 9);
  assign w416[24] = |(datain[215:212] ^ 8);
  assign w416[25] = |(datain[211:208] ^ 1);
  assign w416[26] = |(datain[207:204] ^ 15);
  assign w416[27] = |(datain[203:200] ^ 14);
  assign w416[28] = |(datain[199:196] ^ 11);
  assign w416[29] = |(datain[195:192] ^ 4);
  assign w416[30] = |(datain[191:188] ^ 10);
  assign w416[31] = |(datain[187:184] ^ 3);
  assign w416[32] = |(datain[183:180] ^ 7);
  assign w416[33] = |(datain[179:176] ^ 5);
  assign w416[34] = |(datain[175:172] ^ 0);
  assign w416[35] = |(datain[171:168] ^ 3);
  assign w416[36] = |(datain[167:164] ^ 11);
  assign w416[37] = |(datain[163:160] ^ 15);
  assign w416[38] = |(datain[159:156] ^ 10);
  assign w416[39] = |(datain[155:152] ^ 3);
  assign w416[40] = |(datain[151:148] ^ 10);
  assign w416[41] = |(datain[147:144] ^ 3);
  assign w416[42] = |(datain[143:140] ^ 15);
  assign w416[43] = |(datain[139:136] ^ 11);
  assign comp[416] = ~(|w416);
  wire [74-1:0] w417;
  assign w417[0] = |(datain[311:308] ^ 5);
  assign w417[1] = |(datain[307:304] ^ 11);
  assign w417[2] = |(datain[303:300] ^ 8);
  assign w417[3] = |(datain[299:296] ^ 3);
  assign w417[4] = |(datain[295:292] ^ 14);
  assign w417[5] = |(datain[291:288] ^ 11);
  assign w417[6] = |(datain[287:284] ^ 2);
  assign w417[7] = |(datain[283:280] ^ 0);
  assign w417[8] = |(datain[279:276] ^ 5);
  assign w417[9] = |(datain[275:272] ^ 3);
  assign w417[10] = |(datain[271:268] ^ 11);
  assign w417[11] = |(datain[267:264] ^ 4);
  assign w417[12] = |(datain[263:260] ^ 2);
  assign w417[13] = |(datain[259:256] ^ 10);
  assign w417[14] = |(datain[255:252] ^ 12);
  assign w417[15] = |(datain[251:248] ^ 13);
  assign w417[16] = |(datain[247:244] ^ 2);
  assign w417[17] = |(datain[243:240] ^ 1);
  assign w417[18] = |(datain[239:236] ^ 8);
  assign w417[19] = |(datain[235:232] ^ 0);
  assign w417[20] = |(datain[231:228] ^ 15);
  assign w417[21] = |(datain[227:224] ^ 10);
  assign w417[22] = |(datain[223:220] ^ 0);
  assign w417[23] = |(datain[219:216] ^ 5);
  assign w417[24] = |(datain[215:212] ^ 7);
  assign w417[25] = |(datain[211:208] ^ 5);
  assign w417[26] = |(datain[207:204] ^ 1);
  assign w417[27] = |(datain[203:200] ^ 2);
  assign w417[28] = |(datain[199:196] ^ 8);
  assign w417[29] = |(datain[195:192] ^ 0);
  assign w417[30] = |(datain[191:188] ^ 15);
  assign w417[31] = |(datain[187:184] ^ 14);
  assign w417[32] = |(datain[183:180] ^ 0);
  assign w417[33] = |(datain[179:176] ^ 10);
  assign w417[34] = |(datain[175:172] ^ 7);
  assign w417[35] = |(datain[171:168] ^ 5);
  assign w417[36] = |(datain[167:164] ^ 0);
  assign w417[37] = |(datain[163:160] ^ 13);
  assign w417[38] = |(datain[159:156] ^ 11);
  assign w417[39] = |(datain[155:152] ^ 0);
  assign w417[40] = |(datain[151:148] ^ 0);
  assign w417[41] = |(datain[147:144] ^ 0);
  assign w417[42] = |(datain[143:140] ^ 11);
  assign w417[43] = |(datain[139:136] ^ 9);
  assign w417[44] = |(datain[135:132] ^ 0);
  assign w417[45] = |(datain[131:128] ^ 13);
  assign w417[46] = |(datain[127:124] ^ 0);
  assign w417[47] = |(datain[123:120] ^ 0);
  assign w417[48] = |(datain[119:116] ^ 11);
  assign w417[49] = |(datain[115:112] ^ 10);
  assign w417[50] = |(datain[111:108] ^ 0);
  assign w417[51] = |(datain[107:104] ^ 1);
  assign w417[52] = |(datain[103:100] ^ 0);
  assign w417[53] = |(datain[99:96] ^ 0);
  assign w417[54] = |(datain[95:92] ^ 11);
  assign w417[55] = |(datain[91:88] ^ 11);
  assign w417[56] = |(datain[87:84] ^ 0);
  assign w417[57] = |(datain[83:80] ^ 0);
  assign w417[58] = |(datain[79:76] ^ 0);
  assign w417[59] = |(datain[75:72] ^ 1);
  assign w417[60] = |(datain[71:68] ^ 12);
  assign w417[61] = |(datain[67:64] ^ 13);
  assign w417[62] = |(datain[63:60] ^ 2);
  assign w417[63] = |(datain[59:56] ^ 6);
  assign w417[64] = |(datain[55:52] ^ 11);
  assign w417[65] = |(datain[51:48] ^ 14);
  assign w417[66] = |(datain[47:44] ^ 3);
  assign w417[67] = |(datain[43:40] ^ 4);
  assign w417[68] = |(datain[39:36] ^ 1);
  assign w417[69] = |(datain[35:32] ^ 2);
  assign w417[70] = |(datain[31:28] ^ 11);
  assign w417[71] = |(datain[27:24] ^ 4);
  assign w417[72] = |(datain[23:20] ^ 3);
  assign w417[73] = |(datain[19:16] ^ 0);
  assign comp[417] = ~(|w417);
  wire [40-1:0] w418;
  assign w418[0] = |(datain[311:308] ^ 7);
  assign w418[1] = |(datain[307:304] ^ 5);
  assign w418[2] = |(datain[303:300] ^ 0);
  assign w418[3] = |(datain[299:296] ^ 3);
  assign w418[4] = |(datain[295:292] ^ 14);
  assign w418[5] = |(datain[291:288] ^ 9);
  assign w418[6] = |(datain[287:284] ^ 15);
  assign w418[7] = |(datain[283:280] ^ 8);
  assign w418[8] = |(datain[279:276] ^ 0);
  assign w418[9] = |(datain[275:272] ^ 0);
  assign w418[10] = |(datain[271:268] ^ 8);
  assign w418[11] = |(datain[267:264] ^ 0);
  assign w418[12] = |(datain[263:260] ^ 15);
  assign w418[13] = |(datain[259:256] ^ 12);
  assign w418[14] = |(datain[255:252] ^ 3);
  assign w418[15] = |(datain[251:248] ^ 0);
  assign w418[16] = |(datain[247:244] ^ 7);
  assign w418[17] = |(datain[243:240] ^ 5);
  assign w418[18] = |(datain[239:236] ^ 0);
  assign w418[19] = |(datain[235:232] ^ 9);
  assign w418[20] = |(datain[231:228] ^ 8);
  assign w418[21] = |(datain[227:224] ^ 1);
  assign w418[22] = |(datain[223:220] ^ 15);
  assign w418[23] = |(datain[219:216] ^ 14);
  assign w418[24] = |(datain[215:212] ^ 15);
  assign w418[25] = |(datain[211:208] ^ 13);
  assign w418[26] = |(datain[207:204] ^ 12);
  assign w418[27] = |(datain[203:200] ^ 13);
  assign w418[28] = |(datain[199:196] ^ 7);
  assign w418[29] = |(datain[195:192] ^ 5);
  assign w418[30] = |(datain[191:188] ^ 0);
  assign w418[31] = |(datain[187:184] ^ 3);
  assign w418[32] = |(datain[183:180] ^ 11);
  assign w418[33] = |(datain[179:176] ^ 15);
  assign w418[34] = |(datain[175:172] ^ 12);
  assign w418[35] = |(datain[171:168] ^ 13);
  assign w418[36] = |(datain[167:164] ^ 10);
  assign w418[37] = |(datain[163:160] ^ 11);
  assign w418[38] = |(datain[159:156] ^ 15);
  assign w418[39] = |(datain[155:152] ^ 11);
  assign comp[418] = ~(|w418);
  wire [40-1:0] w419;
  assign w419[0] = |(datain[311:308] ^ 7);
  assign w419[1] = |(datain[307:304] ^ 5);
  assign w419[2] = |(datain[303:300] ^ 0);
  assign w419[3] = |(datain[299:296] ^ 3);
  assign w419[4] = |(datain[295:292] ^ 14);
  assign w419[5] = |(datain[291:288] ^ 9);
  assign w419[6] = |(datain[287:284] ^ 14);
  assign w419[7] = |(datain[283:280] ^ 8);
  assign w419[8] = |(datain[279:276] ^ 0);
  assign w419[9] = |(datain[275:272] ^ 0);
  assign w419[10] = |(datain[271:268] ^ 8);
  assign w419[11] = |(datain[267:264] ^ 0);
  assign w419[12] = |(datain[263:260] ^ 15);
  assign w419[13] = |(datain[259:256] ^ 12);
  assign w419[14] = |(datain[255:252] ^ 3);
  assign w419[15] = |(datain[251:248] ^ 0);
  assign w419[16] = |(datain[247:244] ^ 7);
  assign w419[17] = |(datain[243:240] ^ 5);
  assign w419[18] = |(datain[239:236] ^ 0);
  assign w419[19] = |(datain[235:232] ^ 9);
  assign w419[20] = |(datain[231:228] ^ 8);
  assign w419[21] = |(datain[227:224] ^ 1);
  assign w419[22] = |(datain[223:220] ^ 15);
  assign w419[23] = |(datain[219:216] ^ 14);
  assign w419[24] = |(datain[215:212] ^ 3);
  assign w419[25] = |(datain[211:208] ^ 4);
  assign w419[26] = |(datain[207:204] ^ 1);
  assign w419[27] = |(datain[203:200] ^ 2);
  assign w419[28] = |(datain[199:196] ^ 7);
  assign w419[29] = |(datain[195:192] ^ 5);
  assign w419[30] = |(datain[191:188] ^ 0);
  assign w419[31] = |(datain[187:184] ^ 3);
  assign w419[32] = |(datain[183:180] ^ 11);
  assign w419[33] = |(datain[179:176] ^ 15);
  assign w419[34] = |(datain[175:172] ^ 13);
  assign w419[35] = |(datain[171:168] ^ 13);
  assign w419[36] = |(datain[167:164] ^ 15);
  assign w419[37] = |(datain[163:160] ^ 15);
  assign w419[38] = |(datain[159:156] ^ 15);
  assign w419[39] = |(datain[155:152] ^ 11);
  assign comp[419] = ~(|w419);
  wire [40-1:0] w420;
  assign w420[0] = |(datain[311:308] ^ 7);
  assign w420[1] = |(datain[307:304] ^ 5);
  assign w420[2] = |(datain[303:300] ^ 0);
  assign w420[3] = |(datain[299:296] ^ 3);
  assign w420[4] = |(datain[295:292] ^ 14);
  assign w420[5] = |(datain[291:288] ^ 9);
  assign w420[6] = |(datain[287:284] ^ 4);
  assign w420[7] = |(datain[283:280] ^ 15);
  assign w420[8] = |(datain[279:276] ^ 15);
  assign w420[9] = |(datain[275:272] ^ 14);
  assign w420[10] = |(datain[271:268] ^ 8);
  assign w420[11] = |(datain[267:264] ^ 0);
  assign w420[12] = |(datain[263:260] ^ 15);
  assign w420[13] = |(datain[259:256] ^ 12);
  assign w420[14] = |(datain[255:252] ^ 3);
  assign w420[15] = |(datain[251:248] ^ 0);
  assign w420[16] = |(datain[247:244] ^ 7);
  assign w420[17] = |(datain[243:240] ^ 5);
  assign w420[18] = |(datain[239:236] ^ 0);
  assign w420[19] = |(datain[235:232] ^ 9);
  assign w420[20] = |(datain[231:228] ^ 8);
  assign w420[21] = |(datain[227:224] ^ 1);
  assign w420[22] = |(datain[223:220] ^ 15);
  assign w420[23] = |(datain[219:216] ^ 14);
  assign w420[24] = |(datain[215:212] ^ 15);
  assign w420[25] = |(datain[211:208] ^ 14);
  assign w420[26] = |(datain[207:204] ^ 12);
  assign w420[27] = |(datain[203:200] ^ 13);
  assign w420[28] = |(datain[199:196] ^ 7);
  assign w420[29] = |(datain[195:192] ^ 5);
  assign w420[30] = |(datain[191:188] ^ 0);
  assign w420[31] = |(datain[187:184] ^ 3);
  assign w420[32] = |(datain[183:180] ^ 11);
  assign w420[33] = |(datain[179:176] ^ 15);
  assign w420[34] = |(datain[175:172] ^ 3);
  assign w420[35] = |(datain[171:168] ^ 13);
  assign w420[36] = |(datain[167:164] ^ 1);
  assign w420[37] = |(datain[163:160] ^ 11);
  assign w420[38] = |(datain[159:156] ^ 15);
  assign w420[39] = |(datain[155:152] ^ 11);
  assign comp[420] = ~(|w420);
  wire [44-1:0] w421;
  assign w421[0] = |(datain[311:308] ^ 13);
  assign w421[1] = |(datain[307:304] ^ 15);
  assign w421[2] = |(datain[303:300] ^ 10);
  assign w421[3] = |(datain[299:296] ^ 15);
  assign w421[4] = |(datain[295:292] ^ 11);
  assign w421[5] = |(datain[291:288] ^ 4);
  assign w421[6] = |(datain[287:284] ^ 3);
  assign w421[7] = |(datain[283:280] ^ 0);
  assign w421[8] = |(datain[279:276] ^ 12);
  assign w421[9] = |(datain[275:272] ^ 13);
  assign w421[10] = |(datain[271:268] ^ 2);
  assign w421[11] = |(datain[267:264] ^ 1);
  assign w421[12] = |(datain[263:260] ^ 8);
  assign w421[13] = |(datain[259:256] ^ 1);
  assign w421[14] = |(datain[255:252] ^ 15);
  assign w421[15] = |(datain[251:248] ^ 15);
  assign w421[16] = |(datain[247:244] ^ 12);
  assign w421[17] = |(datain[243:240] ^ 3);
  assign w421[18] = |(datain[239:236] ^ 12);
  assign w421[19] = |(datain[235:232] ^ 3);
  assign w421[20] = |(datain[231:228] ^ 7);
  assign w421[21] = |(datain[227:224] ^ 5);
  assign w421[22] = |(datain[223:220] ^ 1);
  assign w421[23] = |(datain[219:216] ^ 12);
  assign w421[24] = |(datain[215:212] ^ 8);
  assign w421[25] = |(datain[211:208] ^ 12);
  assign w421[26] = |(datain[207:204] ^ 12);
  assign w421[27] = |(datain[203:200] ^ 11);
  assign w421[28] = |(datain[199:196] ^ 2);
  assign w421[29] = |(datain[195:192] ^ 14);
  assign w421[30] = |(datain[191:188] ^ 10);
  assign w421[31] = |(datain[187:184] ^ 1);
  assign w421[32] = |(datain[183:180] ^ 1);
  assign w421[33] = |(datain[179:176] ^ 8);
  assign w421[34] = |(datain[175:172] ^ 0);
  assign w421[35] = |(datain[171:168] ^ 3);
  assign w421[36] = |(datain[167:164] ^ 2);
  assign w421[37] = |(datain[163:160] ^ 11);
  assign w421[38] = |(datain[159:156] ^ 13);
  assign w421[39] = |(datain[155:152] ^ 8);
  assign w421[40] = |(datain[151:148] ^ 2);
  assign w421[41] = |(datain[147:144] ^ 14);
  assign w421[42] = |(datain[143:140] ^ 8);
  assign w421[43] = |(datain[139:136] ^ 9);
  assign comp[421] = ~(|w421);
  wire [42-1:0] w422;
  assign w422[0] = |(datain[311:308] ^ 11);
  assign w422[1] = |(datain[307:304] ^ 4);
  assign w422[2] = |(datain[303:300] ^ 3);
  assign w422[3] = |(datain[299:296] ^ 0);
  assign w422[4] = |(datain[295:292] ^ 12);
  assign w422[5] = |(datain[291:288] ^ 13);
  assign w422[6] = |(datain[287:284] ^ 2);
  assign w422[7] = |(datain[283:280] ^ 1);
  assign w422[8] = |(datain[279:276] ^ 8);
  assign w422[9] = |(datain[275:272] ^ 1);
  assign w422[10] = |(datain[271:268] ^ 15);
  assign w422[11] = |(datain[267:264] ^ 15);
  assign w422[12] = |(datain[263:260] ^ 3);
  assign w422[13] = |(datain[259:256] ^ 13);
  assign w422[14] = |(datain[255:252] ^ 1);
  assign w422[15] = |(datain[251:248] ^ 11);
  assign w422[16] = |(datain[247:244] ^ 7);
  assign w422[17] = |(datain[243:240] ^ 5);
  assign w422[18] = |(datain[239:236] ^ 1);
  assign w422[19] = |(datain[235:232] ^ 7);
  assign w422[20] = |(datain[231:228] ^ 11);
  assign w422[21] = |(datain[227:224] ^ 14);
  assign w422[22] = |(datain[223:220] ^ 1);
  assign w422[23] = |(datain[219:216] ^ 11);
  assign w422[24] = |(datain[215:212] ^ 0);
  assign w422[25] = |(datain[211:208] ^ 4);
  assign w422[26] = |(datain[207:204] ^ 5);
  assign w422[27] = |(datain[203:200] ^ 11);
  assign w422[28] = |(datain[199:196] ^ 8);
  assign w422[29] = |(datain[195:192] ^ 1);
  assign w422[30] = |(datain[191:188] ^ 14);
  assign w422[31] = |(datain[187:184] ^ 11);
  assign w422[32] = |(datain[183:180] ^ 0);
  assign w422[33] = |(datain[179:176] ^ 0);
  assign w422[34] = |(datain[175:172] ^ 0);
  assign w422[35] = |(datain[171:168] ^ 1);
  assign w422[36] = |(datain[167:164] ^ 0);
  assign w422[37] = |(datain[163:160] ^ 3);
  assign w422[38] = |(datain[159:156] ^ 15);
  assign w422[39] = |(datain[155:152] ^ 3);
  assign w422[40] = |(datain[151:148] ^ 11);
  assign w422[41] = |(datain[147:144] ^ 15);
  assign comp[422] = ~(|w422);
  wire [34-1:0] w423;
  assign w423[0] = |(datain[311:308] ^ 5);
  assign w423[1] = |(datain[307:304] ^ 0);
  assign w423[2] = |(datain[303:300] ^ 14);
  assign w423[3] = |(datain[299:296] ^ 8);
  assign w423[4] = |(datain[295:292] ^ 0);
  assign w423[5] = |(datain[291:288] ^ 0);
  assign w423[6] = |(datain[287:284] ^ 0);
  assign w423[7] = |(datain[283:280] ^ 0);
  assign w423[8] = |(datain[279:276] ^ 5);
  assign w423[9] = |(datain[275:272] ^ 14);
  assign w423[10] = |(datain[271:268] ^ 8);
  assign w423[11] = |(datain[267:264] ^ 3);
  assign w423[12] = |(datain[263:260] ^ 12);
  assign w423[13] = |(datain[259:256] ^ 6);
  assign w423[14] = |(datain[255:252] ^ 0);
  assign w423[15] = |(datain[251:248] ^ 13);
  assign w423[16] = |(datain[247:244] ^ 11);
  assign w423[17] = |(datain[243:240] ^ 9);
  assign w423[18] = |(datain[239:236] ^ 2);
  assign w423[19] = |(datain[235:232] ^ 5);
  assign w423[20] = |(datain[231:228] ^ 0);
  assign w423[21] = |(datain[227:224] ^ 0);
  assign w423[22] = |(datain[223:220] ^ 3);
  assign w423[23] = |(datain[219:216] ^ 1);
  assign w423[24] = |(datain[215:212] ^ 0);
  assign w423[25] = |(datain[211:208] ^ 12);
  assign w423[26] = |(datain[207:204] ^ 4);
  assign w423[27] = |(datain[203:200] ^ 6);
  assign w423[28] = |(datain[199:196] ^ 4);
  assign w423[29] = |(datain[195:192] ^ 9);
  assign w423[30] = |(datain[191:188] ^ 7);
  assign w423[31] = |(datain[187:184] ^ 5);
  assign w423[32] = |(datain[183:180] ^ 15);
  assign w423[33] = |(datain[179:176] ^ 10);
  assign comp[423] = ~(|w423);
  wire [74-1:0] w424;
  assign w424[0] = |(datain[311:308] ^ 11);
  assign w424[1] = |(datain[307:304] ^ 9);
  assign w424[2] = |(datain[303:300] ^ 0);
  assign w424[3] = |(datain[299:296] ^ 3);
  assign w424[4] = |(datain[295:292] ^ 0);
  assign w424[5] = |(datain[291:288] ^ 0);
  assign w424[6] = |(datain[287:284] ^ 11);
  assign w424[7] = |(datain[283:280] ^ 4);
  assign w424[8] = |(datain[279:276] ^ 4);
  assign w424[9] = |(datain[275:272] ^ 0);
  assign w424[10] = |(datain[271:268] ^ 12);
  assign w424[11] = |(datain[267:264] ^ 13);
  assign w424[12] = |(datain[263:260] ^ 2);
  assign w424[13] = |(datain[259:256] ^ 1);
  assign w424[14] = |(datain[255:252] ^ 2);
  assign w424[15] = |(datain[251:248] ^ 14);
  assign w424[16] = |(datain[247:244] ^ 8);
  assign w424[17] = |(datain[243:240] ^ 11);
  assign w424[18] = |(datain[239:236] ^ 1);
  assign w424[19] = |(datain[235:232] ^ 14);
  assign w424[20] = |(datain[231:228] ^ 10);
  assign w424[21] = |(datain[227:224] ^ 4);
  assign w424[22] = |(datain[223:220] ^ 0);
  assign w424[23] = |(datain[219:216] ^ 2);
  assign w424[24] = |(datain[215:212] ^ 5);
  assign w424[25] = |(datain[211:208] ^ 3);
  assign w424[26] = |(datain[207:204] ^ 11);
  assign w424[27] = |(datain[203:200] ^ 0);
  assign w424[28] = |(datain[199:196] ^ 0);
  assign w424[29] = |(datain[195:192] ^ 2);
  assign w424[30] = |(datain[191:188] ^ 3);
  assign w424[31] = |(datain[187:184] ^ 3);
  assign w424[32] = |(datain[183:180] ^ 12);
  assign w424[33] = |(datain[179:176] ^ 9);
  assign w424[34] = |(datain[175:172] ^ 3);
  assign w424[35] = |(datain[171:168] ^ 3);
  assign w424[36] = |(datain[167:164] ^ 13);
  assign w424[37] = |(datain[163:160] ^ 2);
  assign w424[38] = |(datain[159:156] ^ 11);
  assign w424[39] = |(datain[155:152] ^ 4);
  assign w424[40] = |(datain[151:148] ^ 4);
  assign w424[41] = |(datain[147:144] ^ 2);
  assign w424[42] = |(datain[143:140] ^ 12);
  assign w424[43] = |(datain[139:136] ^ 13);
  assign w424[44] = |(datain[135:132] ^ 2);
  assign w424[45] = |(datain[131:128] ^ 1);
  assign w424[46] = |(datain[127:124] ^ 2);
  assign w424[47] = |(datain[123:120] ^ 14);
  assign w424[48] = |(datain[119:116] ^ 8);
  assign w424[49] = |(datain[115:112] ^ 14);
  assign w424[50] = |(datain[111:108] ^ 1);
  assign w424[51] = |(datain[107:104] ^ 14);
  assign w424[52] = |(datain[103:100] ^ 11);
  assign w424[53] = |(datain[99:96] ^ 9);
  assign w424[54] = |(datain[95:92] ^ 0);
  assign w424[55] = |(datain[91:88] ^ 2);
  assign w424[56] = |(datain[87:84] ^ 3);
  assign w424[57] = |(datain[83:80] ^ 3);
  assign w424[58] = |(datain[79:76] ^ 13);
  assign w424[59] = |(datain[75:72] ^ 2);
  assign w424[60] = |(datain[71:68] ^ 5);
  assign w424[61] = |(datain[67:64] ^ 11);
  assign w424[62] = |(datain[63:60] ^ 11);
  assign w424[63] = |(datain[59:56] ^ 9);
  assign w424[64] = |(datain[55:52] ^ 15);
  assign w424[65] = |(datain[51:48] ^ 8);
  assign w424[66] = |(datain[47:44] ^ 0);
  assign w424[67] = |(datain[43:40] ^ 3);
  assign w424[68] = |(datain[39:36] ^ 11);
  assign w424[69] = |(datain[35:32] ^ 4);
  assign w424[70] = |(datain[31:28] ^ 4);
  assign w424[71] = |(datain[27:24] ^ 0);
  assign w424[72] = |(datain[23:20] ^ 12);
  assign w424[73] = |(datain[19:16] ^ 13);
  assign comp[424] = ~(|w424);
  wire [74-1:0] w425;
  assign w425[0] = |(datain[311:308] ^ 12);
  assign w425[1] = |(datain[307:304] ^ 5);
  assign w425[2] = |(datain[303:300] ^ 0);
  assign w425[3] = |(datain[299:296] ^ 2);
  assign w425[4] = |(datain[295:292] ^ 11);
  assign w425[5] = |(datain[291:288] ^ 9);
  assign w425[6] = |(datain[287:284] ^ 0);
  assign w425[7] = |(datain[283:280] ^ 3);
  assign w425[8] = |(datain[279:276] ^ 0);
  assign w425[9] = |(datain[275:272] ^ 0);
  assign w425[10] = |(datain[271:268] ^ 11);
  assign w425[11] = |(datain[267:264] ^ 4);
  assign w425[12] = |(datain[263:260] ^ 4);
  assign w425[13] = |(datain[259:256] ^ 0);
  assign w425[14] = |(datain[255:252] ^ 12);
  assign w425[15] = |(datain[251:248] ^ 13);
  assign w425[16] = |(datain[247:244] ^ 2);
  assign w425[17] = |(datain[243:240] ^ 1);
  assign w425[18] = |(datain[239:236] ^ 2);
  assign w425[19] = |(datain[235:232] ^ 14);
  assign w425[20] = |(datain[231:228] ^ 8);
  assign w425[21] = |(datain[227:224] ^ 11);
  assign w425[22] = |(datain[223:220] ^ 1);
  assign w425[23] = |(datain[219:216] ^ 14);
  assign w425[24] = |(datain[215:212] ^ 12);
  assign w425[25] = |(datain[211:208] ^ 1);
  assign w425[26] = |(datain[207:204] ^ 0);
  assign w425[27] = |(datain[203:200] ^ 2);
  assign w425[28] = |(datain[199:196] ^ 5);
  assign w425[29] = |(datain[195:192] ^ 3);
  assign w425[30] = |(datain[191:188] ^ 11);
  assign w425[31] = |(datain[187:184] ^ 0);
  assign w425[32] = |(datain[183:180] ^ 0);
  assign w425[33] = |(datain[179:176] ^ 2);
  assign w425[34] = |(datain[175:172] ^ 3);
  assign w425[35] = |(datain[171:168] ^ 3);
  assign w425[36] = |(datain[167:164] ^ 12);
  assign w425[37] = |(datain[163:160] ^ 9);
  assign w425[38] = |(datain[159:156] ^ 3);
  assign w425[39] = |(datain[155:152] ^ 3);
  assign w425[40] = |(datain[151:148] ^ 13);
  assign w425[41] = |(datain[147:144] ^ 2);
  assign w425[42] = |(datain[143:140] ^ 11);
  assign w425[43] = |(datain[139:136] ^ 4);
  assign w425[44] = |(datain[135:132] ^ 4);
  assign w425[45] = |(datain[131:128] ^ 2);
  assign w425[46] = |(datain[127:124] ^ 12);
  assign w425[47] = |(datain[123:120] ^ 13);
  assign w425[48] = |(datain[119:116] ^ 2);
  assign w425[49] = |(datain[115:112] ^ 1);
  assign w425[50] = |(datain[111:108] ^ 2);
  assign w425[51] = |(datain[107:104] ^ 14);
  assign w425[52] = |(datain[103:100] ^ 8);
  assign w425[53] = |(datain[99:96] ^ 14);
  assign w425[54] = |(datain[95:92] ^ 1);
  assign w425[55] = |(datain[91:88] ^ 14);
  assign w425[56] = |(datain[87:84] ^ 13);
  assign w425[57] = |(datain[83:80] ^ 6);
  assign w425[58] = |(datain[79:76] ^ 0);
  assign w425[59] = |(datain[75:72] ^ 2);
  assign w425[60] = |(datain[71:68] ^ 3);
  assign w425[61] = |(datain[67:64] ^ 3);
  assign w425[62] = |(datain[63:60] ^ 13);
  assign w425[63] = |(datain[59:56] ^ 2);
  assign w425[64] = |(datain[55:52] ^ 5);
  assign w425[65] = |(datain[51:48] ^ 11);
  assign w425[66] = |(datain[47:44] ^ 11);
  assign w425[67] = |(datain[43:40] ^ 9);
  assign w425[68] = |(datain[39:36] ^ 14);
  assign w425[69] = |(datain[35:32] ^ 6);
  assign w425[70] = |(datain[31:28] ^ 0);
  assign w425[71] = |(datain[27:24] ^ 3);
  assign w425[72] = |(datain[23:20] ^ 11);
  assign w425[73] = |(datain[19:16] ^ 4);
  assign comp[425] = ~(|w425);
  wire [44-1:0] w426;
  assign w426[0] = |(datain[311:308] ^ 8);
  assign w426[1] = |(datain[307:304] ^ 13);
  assign w426[2] = |(datain[303:300] ^ 5);
  assign w426[3] = |(datain[299:296] ^ 6);
  assign w426[4] = |(datain[295:292] ^ 8);
  assign w426[5] = |(datain[291:288] ^ 8);
  assign w426[6] = |(datain[287:284] ^ 9);
  assign w426[7] = |(datain[283:280] ^ 0);
  assign w426[8] = |(datain[279:276] ^ 11);
  assign w426[9] = |(datain[275:272] ^ 9);
  assign w426[10] = |(datain[271:268] ^ 3);
  assign w426[11] = |(datain[267:264] ^ 15);
  assign w426[12] = |(datain[263:260] ^ 0);
  assign w426[13] = |(datain[259:256] ^ 0);
  assign w426[14] = |(datain[255:252] ^ 12);
  assign w426[15] = |(datain[251:248] ^ 13);
  assign w426[16] = |(datain[247:244] ^ 2);
  assign w426[17] = |(datain[243:240] ^ 1);
  assign w426[18] = |(datain[239:236] ^ 7);
  assign w426[19] = |(datain[235:232] ^ 2);
  assign w426[20] = |(datain[231:228] ^ 1);
  assign w426[21] = |(datain[227:224] ^ 10);
  assign w426[22] = |(datain[223:220] ^ 8);
  assign w426[23] = |(datain[219:216] ^ 13);
  assign w426[24] = |(datain[215:212] ^ 9);
  assign w426[25] = |(datain[211:208] ^ 6);
  assign w426[26] = |(datain[207:204] ^ 12);
  assign w426[27] = |(datain[203:200] ^ 13);
  assign w426[28] = |(datain[199:196] ^ 0);
  assign w426[29] = |(datain[195:192] ^ 0);
  assign w426[30] = |(datain[191:188] ^ 11);
  assign w426[31] = |(datain[187:184] ^ 8);
  assign w426[32] = |(datain[183:180] ^ 0);
  assign w426[33] = |(datain[179:176] ^ 2);
  assign w426[34] = |(datain[175:172] ^ 3);
  assign w426[35] = |(datain[171:168] ^ 13);
  assign w426[36] = |(datain[167:164] ^ 12);
  assign w426[37] = |(datain[163:160] ^ 13);
  assign w426[38] = |(datain[159:156] ^ 2);
  assign w426[39] = |(datain[155:152] ^ 1);
  assign w426[40] = |(datain[151:148] ^ 7);
  assign w426[41] = |(datain[147:144] ^ 2);
  assign w426[42] = |(datain[143:140] ^ 0);
  assign w426[43] = |(datain[139:136] ^ 9);
  assign comp[426] = ~(|w426);
  wire [70-1:0] w427;
  assign w427[0] = |(datain[311:308] ^ 12);
  assign w427[1] = |(datain[307:304] ^ 3);
  assign w427[2] = |(datain[303:300] ^ 5);
  assign w427[3] = |(datain[299:296] ^ 3);
  assign w427[4] = |(datain[295:292] ^ 8);
  assign w427[5] = |(datain[291:288] ^ 11);
  assign w427[6] = |(datain[287:284] ^ 9);
  assign w427[7] = |(datain[283:280] ^ 15);
  assign w427[8] = |(datain[279:276] ^ 0);
  assign w427[9] = |(datain[275:272] ^ 4);
  assign w427[10] = |(datain[271:268] ^ 1);
  assign w427[11] = |(datain[267:264] ^ 0);
  assign w427[12] = |(datain[263:260] ^ 12);
  assign w427[13] = |(datain[259:256] ^ 13);
  assign w427[14] = |(datain[255:252] ^ 2);
  assign w427[15] = |(datain[251:248] ^ 1);
  assign w427[16] = |(datain[247:244] ^ 5);
  assign w427[17] = |(datain[243:240] ^ 11);
  assign w427[18] = |(datain[239:236] ^ 12);
  assign w427[19] = |(datain[235:232] ^ 3);
  assign w427[20] = |(datain[231:228] ^ 11);
  assign w427[21] = |(datain[227:224] ^ 4);
  assign w427[22] = |(datain[223:220] ^ 3);
  assign w427[23] = |(datain[219:216] ^ 15);
  assign w427[24] = |(datain[215:212] ^ 14);
  assign w427[25] = |(datain[211:208] ^ 8);
  assign w427[26] = |(datain[207:204] ^ 15);
  assign w427[27] = |(datain[203:200] ^ 2);
  assign w427[28] = |(datain[199:196] ^ 15);
  assign w427[29] = |(datain[195:192] ^ 15);
  assign w427[30] = |(datain[191:188] ^ 12);
  assign w427[31] = |(datain[187:184] ^ 3);
  assign w427[32] = |(datain[183:180] ^ 11);
  assign w427[33] = |(datain[179:176] ^ 4);
  assign w427[34] = |(datain[175:172] ^ 4);
  assign w427[35] = |(datain[171:168] ^ 0);
  assign w427[36] = |(datain[167:164] ^ 14);
  assign w427[37] = |(datain[163:160] ^ 8);
  assign w427[38] = |(datain[159:156] ^ 14);
  assign w427[39] = |(datain[155:152] ^ 12);
  assign w427[40] = |(datain[151:148] ^ 15);
  assign w427[41] = |(datain[147:144] ^ 15);
  assign w427[42] = |(datain[143:140] ^ 12);
  assign w427[43] = |(datain[139:136] ^ 3);
  assign w427[44] = |(datain[135:132] ^ 11);
  assign w427[45] = |(datain[131:128] ^ 4);
  assign w427[46] = |(datain[127:124] ^ 4);
  assign w427[47] = |(datain[123:120] ^ 3);
  assign w427[48] = |(datain[119:116] ^ 8);
  assign w427[49] = |(datain[115:112] ^ 11);
  assign w427[50] = |(datain[111:108] ^ 13);
  assign w427[51] = |(datain[107:104] ^ 3);
  assign w427[52] = |(datain[103:100] ^ 8);
  assign w427[53] = |(datain[99:96] ^ 1);
  assign w427[54] = |(datain[95:92] ^ 12);
  assign w427[55] = |(datain[91:88] ^ 2);
  assign w427[56] = |(datain[87:84] ^ 1);
  assign w427[57] = |(datain[83:80] ^ 14);
  assign w427[58] = |(datain[79:76] ^ 0);
  assign w427[59] = |(datain[75:72] ^ 4);
  assign w427[60] = |(datain[71:68] ^ 12);
  assign w427[61] = |(datain[67:64] ^ 13);
  assign w427[62] = |(datain[63:60] ^ 2);
  assign w427[63] = |(datain[59:56] ^ 1);
  assign w427[64] = |(datain[55:52] ^ 12);
  assign w427[65] = |(datain[51:48] ^ 3);
  assign w427[66] = |(datain[47:44] ^ 11);
  assign w427[67] = |(datain[43:40] ^ 4);
  assign w427[68] = |(datain[39:36] ^ 2);
  assign w427[69] = |(datain[35:32] ^ 10);
  assign comp[427] = ~(|w427);
  wire [42-1:0] w428;
  assign w428[0] = |(datain[311:308] ^ 2);
  assign w428[1] = |(datain[307:304] ^ 3);
  assign w428[2] = |(datain[303:300] ^ 11);
  assign w428[3] = |(datain[299:296] ^ 11);
  assign w428[4] = |(datain[295:292] ^ 2);
  assign w428[5] = |(datain[291:288] ^ 0);
  assign w428[6] = |(datain[287:284] ^ 2);
  assign w428[7] = |(datain[283:280] ^ 8);
  assign w428[8] = |(datain[279:276] ^ 2);
  assign w428[9] = |(datain[275:272] ^ 14);
  assign w428[10] = |(datain[271:268] ^ 0);
  assign w428[11] = |(datain[267:264] ^ 0);
  assign w428[12] = |(datain[263:260] ^ 2);
  assign w428[13] = |(datain[259:256] ^ 7);
  assign w428[14] = |(datain[255:252] ^ 2);
  assign w428[15] = |(datain[251:248] ^ 14);
  assign w428[16] = |(datain[247:244] ^ 3);
  assign w428[17] = |(datain[243:240] ^ 2);
  assign w428[18] = |(datain[239:236] ^ 2);
  assign w428[19] = |(datain[235:232] ^ 7);
  assign w428[20] = |(datain[231:228] ^ 4);
  assign w428[21] = |(datain[227:224] ^ 3);
  assign w428[22] = |(datain[223:220] ^ 8);
  assign w428[23] = |(datain[219:216] ^ 1);
  assign w428[24] = |(datain[215:212] ^ 15);
  assign w428[25] = |(datain[211:208] ^ 11);
  assign w428[26] = |(datain[207:204] ^ 1);
  assign w428[27] = |(datain[203:200] ^ 11);
  assign w428[28] = |(datain[199:196] ^ 2);
  assign w428[29] = |(datain[195:192] ^ 14);
  assign w428[30] = |(datain[191:188] ^ 7);
  assign w428[31] = |(datain[187:184] ^ 5);
  assign w428[32] = |(datain[183:180] ^ 15);
  assign w428[33] = |(datain[179:176] ^ 3);
  assign w428[34] = |(datain[175:172] ^ 14);
  assign w428[35] = |(datain[171:168] ^ 9);
  assign w428[36] = |(datain[167:164] ^ 14);
  assign w428[37] = |(datain[163:160] ^ 13);
  assign w428[38] = |(datain[159:156] ^ 15);
  assign w428[39] = |(datain[155:152] ^ 14);
  assign w428[40] = |(datain[151:148] ^ 14);
  assign w428[41] = |(datain[147:144] ^ 10);
  assign comp[428] = ~(|w428);
  wire [42-1:0] w429;
  assign w429[0] = |(datain[311:308] ^ 8);
  assign w429[1] = |(datain[307:304] ^ 14);
  assign w429[2] = |(datain[303:300] ^ 13);
  assign w429[3] = |(datain[299:296] ^ 10);
  assign w429[4] = |(datain[295:292] ^ 10);
  assign w429[5] = |(datain[291:288] ^ 1);
  assign w429[6] = |(datain[287:284] ^ 0);
  assign w429[7] = |(datain[283:280] ^ 6);
  assign w429[8] = |(datain[279:276] ^ 0);
  assign w429[9] = |(datain[275:272] ^ 0);
  assign w429[10] = |(datain[271:268] ^ 8);
  assign w429[11] = |(datain[267:264] ^ 14);
  assign w429[12] = |(datain[263:260] ^ 13);
  assign w429[13] = |(datain[259:256] ^ 8);
  assign w429[14] = |(datain[255:252] ^ 11);
  assign w429[15] = |(datain[251:248] ^ 9);
  assign w429[16] = |(datain[247:244] ^ 15);
  assign w429[17] = |(datain[243:240] ^ 15);
  assign w429[18] = |(datain[239:236] ^ 15);
  assign w429[19] = |(datain[235:232] ^ 15);
  assign w429[20] = |(datain[231:228] ^ 8);
  assign w429[21] = |(datain[227:224] ^ 11);
  assign w429[22] = |(datain[223:220] ^ 15);
  assign w429[23] = |(datain[219:216] ^ 2);
  assign w429[24] = |(datain[215:212] ^ 8);
  assign w429[25] = |(datain[211:208] ^ 1);
  assign w429[26] = |(datain[207:204] ^ 3);
  assign w429[27] = |(datain[203:200] ^ 12);
  assign w429[28] = |(datain[199:196] ^ 15);
  assign w429[29] = |(datain[195:192] ^ 3);
  assign w429[30] = |(datain[191:188] ^ 10);
  assign w429[31] = |(datain[187:184] ^ 5);
  assign w429[32] = |(datain[183:180] ^ 7);
  assign w429[33] = |(datain[179:176] ^ 4);
  assign w429[34] = |(datain[175:172] ^ 0);
  assign w429[35] = |(datain[171:168] ^ 6);
  assign w429[36] = |(datain[167:164] ^ 4);
  assign w429[37] = |(datain[163:160] ^ 6);
  assign w429[38] = |(datain[159:156] ^ 14);
  assign w429[39] = |(datain[155:152] ^ 2);
  assign w429[40] = |(datain[151:148] ^ 15);
  assign w429[41] = |(datain[147:144] ^ 7);
  assign comp[429] = ~(|w429);
  wire [64-1:0] w430;
  assign w430[0] = |(datain[311:308] ^ 15);
  assign w430[1] = |(datain[307:304] ^ 9);
  assign w430[2] = |(datain[303:300] ^ 0);
  assign w430[3] = |(datain[299:296] ^ 1);
  assign w430[4] = |(datain[295:292] ^ 7);
  assign w430[5] = |(datain[291:288] ^ 5);
  assign w430[6] = |(datain[287:284] ^ 0);
  assign w430[7] = |(datain[283:280] ^ 5);
  assign w430[8] = |(datain[279:276] ^ 8);
  assign w430[9] = |(datain[275:272] ^ 0);
  assign w430[10] = |(datain[271:268] ^ 15);
  assign w430[11] = |(datain[267:264] ^ 12);
  assign w430[12] = |(datain[263:260] ^ 0);
  assign w430[13] = |(datain[259:256] ^ 2);
  assign w430[14] = |(datain[255:252] ^ 7);
  assign w430[15] = |(datain[251:248] ^ 4);
  assign w430[16] = |(datain[247:244] ^ 0);
  assign w430[17] = |(datain[243:240] ^ 3);
  assign w430[18] = |(datain[239:236] ^ 14);
  assign w430[19] = |(datain[235:232] ^ 9);
  assign w430[20] = |(datain[231:228] ^ 9);
  assign w430[21] = |(datain[227:224] ^ 5);
  assign w430[22] = |(datain[223:220] ^ 0);
  assign w430[23] = |(datain[219:216] ^ 0);
  assign w430[24] = |(datain[215:212] ^ 9);
  assign w430[25] = |(datain[211:208] ^ 12);
  assign w430[26] = |(datain[207:204] ^ 2);
  assign w430[27] = |(datain[203:200] ^ 14);
  assign w430[28] = |(datain[199:196] ^ 15);
  assign w430[29] = |(datain[195:192] ^ 15);
  assign w430[30] = |(datain[191:188] ^ 1);
  assign w430[31] = |(datain[187:184] ^ 14);
  assign w430[32] = |(datain[183:180] ^ 8);
  assign w430[33] = |(datain[179:176] ^ 4);
  assign w430[34] = |(datain[175:172] ^ 0);
  assign w430[35] = |(datain[171:168] ^ 1);
  assign w430[36] = |(datain[167:164] ^ 7);
  assign w430[37] = |(datain[163:160] ^ 3);
  assign w430[38] = |(datain[159:156] ^ 0);
  assign w430[39] = |(datain[155:152] ^ 3);
  assign w430[40] = |(datain[151:148] ^ 14);
  assign w430[41] = |(datain[147:144] ^ 9);
  assign w430[42] = |(datain[143:140] ^ 10);
  assign w430[43] = |(datain[139:136] ^ 7);
  assign w430[44] = |(datain[135:132] ^ 0);
  assign w430[45] = |(datain[131:128] ^ 0);
  assign w430[46] = |(datain[127:124] ^ 2);
  assign w430[47] = |(datain[123:120] ^ 6);
  assign w430[48] = |(datain[119:116] ^ 8);
  assign w430[49] = |(datain[115:112] ^ 1);
  assign w430[50] = |(datain[111:108] ^ 11);
  assign w430[51] = |(datain[107:104] ^ 15);
  assign w430[52] = |(datain[103:100] ^ 15);
  assign w430[53] = |(datain[99:96] ^ 0);
  assign w430[54] = |(datain[95:92] ^ 0);
  assign w430[55] = |(datain[91:88] ^ 0);
  assign w430[56] = |(datain[87:84] ^ 8);
  assign w430[57] = |(datain[83:80] ^ 1);
  assign w430[58] = |(datain[79:76] ^ 12);
  assign w430[59] = |(datain[75:72] ^ 6);
  assign w430[60] = |(datain[71:68] ^ 7);
  assign w430[61] = |(datain[67:64] ^ 5);
  assign w430[62] = |(datain[63:60] ^ 0);
  assign w430[63] = |(datain[59:56] ^ 3);
  assign comp[430] = ~(|w430);
  wire [76-1:0] w431;
  assign w431[0] = |(datain[311:308] ^ 0);
  assign w431[1] = |(datain[307:304] ^ 1);
  assign w431[2] = |(datain[303:300] ^ 11);
  assign w431[3] = |(datain[299:296] ^ 4);
  assign w431[4] = |(datain[295:292] ^ 4);
  assign w431[5] = |(datain[291:288] ^ 0);
  assign w431[6] = |(datain[287:284] ^ 12);
  assign w431[7] = |(datain[283:280] ^ 13);
  assign w431[8] = |(datain[279:276] ^ 2);
  assign w431[9] = |(datain[275:272] ^ 1);
  assign w431[10] = |(datain[271:268] ^ 8);
  assign w431[11] = |(datain[267:264] ^ 1);
  assign w431[12] = |(datain[263:260] ^ 12);
  assign w431[13] = |(datain[259:256] ^ 7);
  assign w431[14] = |(datain[255:252] ^ 0);
  assign w431[15] = |(datain[251:248] ^ 0);
  assign w431[16] = |(datain[247:244] ^ 0);
  assign w431[17] = |(datain[243:240] ^ 1);
  assign w431[18] = |(datain[239:236] ^ 8);
  assign w431[19] = |(datain[235:232] ^ 9);
  assign w431[20] = |(datain[231:228] ^ 3);
  assign w431[21] = |(datain[227:224] ^ 14);
  assign w431[22] = |(datain[223:220] ^ 8);
  assign w431[23] = |(datain[219:216] ^ 10);
  assign w431[24] = |(datain[215:212] ^ 0);
  assign w431[25] = |(datain[211:208] ^ 1);
  assign w431[26] = |(datain[207:204] ^ 12);
  assign w431[27] = |(datain[203:200] ^ 6);
  assign w431[28] = |(datain[199:196] ^ 0);
  assign w431[29] = |(datain[195:192] ^ 6);
  assign w431[30] = |(datain[191:188] ^ 8);
  assign w431[31] = |(datain[187:184] ^ 14);
  assign w431[32] = |(datain[183:180] ^ 0);
  assign w431[33] = |(datain[179:176] ^ 1);
  assign w431[34] = |(datain[175:172] ^ 13);
  assign w431[35] = |(datain[171:168] ^ 14);
  assign w431[36] = |(datain[167:164] ^ 11);
  assign w431[37] = |(datain[163:160] ^ 8);
  assign w431[38] = |(datain[159:156] ^ 0);
  assign w431[39] = |(datain[155:152] ^ 0);
  assign w431[40] = |(datain[151:148] ^ 4);
  assign w431[41] = |(datain[147:144] ^ 2);
  assign w431[42] = |(datain[143:140] ^ 3);
  assign w431[43] = |(datain[139:136] ^ 3);
  assign w431[44] = |(datain[135:132] ^ 12);
  assign w431[45] = |(datain[131:128] ^ 9);
  assign w431[46] = |(datain[127:124] ^ 3);
  assign w431[47] = |(datain[123:120] ^ 3);
  assign w431[48] = |(datain[119:116] ^ 13);
  assign w431[49] = |(datain[115:112] ^ 2);
  assign w431[50] = |(datain[111:108] ^ 12);
  assign w431[51] = |(datain[107:104] ^ 13);
  assign w431[52] = |(datain[103:100] ^ 2);
  assign w431[53] = |(datain[99:96] ^ 1);
  assign w431[54] = |(datain[95:92] ^ 11);
  assign w431[55] = |(datain[91:88] ^ 9);
  assign w431[56] = |(datain[87:84] ^ 0);
  assign w431[57] = |(datain[83:80] ^ 6);
  assign w431[58] = |(datain[79:76] ^ 0);
  assign w431[59] = |(datain[75:72] ^ 0);
  assign w431[60] = |(datain[71:68] ^ 11);
  assign w431[61] = |(datain[67:64] ^ 10);
  assign w431[62] = |(datain[63:60] ^ 8);
  assign w431[63] = |(datain[59:56] ^ 9);
  assign w431[64] = |(datain[55:52] ^ 0);
  assign w431[65] = |(datain[51:48] ^ 1);
  assign w431[66] = |(datain[47:44] ^ 11);
  assign w431[67] = |(datain[43:40] ^ 4);
  assign w431[68] = |(datain[39:36] ^ 4);
  assign w431[69] = |(datain[35:32] ^ 0);
  assign w431[70] = |(datain[31:28] ^ 12);
  assign w431[71] = |(datain[27:24] ^ 13);
  assign w431[72] = |(datain[23:20] ^ 2);
  assign w431[73] = |(datain[19:16] ^ 1);
  assign w431[74] = |(datain[15:12] ^ 11);
  assign w431[75] = |(datain[11:8] ^ 4);
  assign comp[431] = ~(|w431);
  wire [74-1:0] w432;
  assign w432[0] = |(datain[311:308] ^ 11);
  assign w432[1] = |(datain[307:304] ^ 9);
  assign w432[2] = |(datain[303:300] ^ 9);
  assign w432[3] = |(datain[299:296] ^ 4);
  assign w432[4] = |(datain[295:292] ^ 0);
  assign w432[5] = |(datain[291:288] ^ 4);
  assign w432[6] = |(datain[287:284] ^ 11);
  assign w432[7] = |(datain[283:280] ^ 10);
  assign w432[8] = |(datain[279:276] ^ 0);
  assign w432[9] = |(datain[275:272] ^ 0);
  assign w432[10] = |(datain[271:268] ^ 0);
  assign w432[11] = |(datain[267:264] ^ 1);
  assign w432[12] = |(datain[263:260] ^ 11);
  assign w432[13] = |(datain[259:256] ^ 4);
  assign w432[14] = |(datain[255:252] ^ 4);
  assign w432[15] = |(datain[251:248] ^ 0);
  assign w432[16] = |(datain[247:244] ^ 14);
  assign w432[17] = |(datain[243:240] ^ 8);
  assign w432[18] = |(datain[239:236] ^ 5);
  assign w432[19] = |(datain[235:232] ^ 4);
  assign w432[20] = |(datain[231:228] ^ 0);
  assign w432[21] = |(datain[227:224] ^ 0);
  assign w432[22] = |(datain[223:220] ^ 7);
  assign w432[23] = |(datain[219:216] ^ 2);
  assign w432[24] = |(datain[215:212] ^ 2);
  assign w432[25] = |(datain[211:208] ^ 6);
  assign w432[26] = |(datain[207:204] ^ 3);
  assign w432[27] = |(datain[203:200] ^ 3);
  assign w432[28] = |(datain[199:196] ^ 13);
  assign w432[29] = |(datain[195:192] ^ 2);
  assign w432[30] = |(datain[191:188] ^ 3);
  assign w432[31] = |(datain[187:184] ^ 3);
  assign w432[32] = |(datain[183:180] ^ 12);
  assign w432[33] = |(datain[179:176] ^ 9);
  assign w432[34] = |(datain[175:172] ^ 11);
  assign w432[35] = |(datain[171:168] ^ 8);
  assign w432[36] = |(datain[167:164] ^ 0);
  assign w432[37] = |(datain[163:160] ^ 0);
  assign w432[38] = |(datain[159:156] ^ 4);
  assign w432[39] = |(datain[155:152] ^ 2);
  assign w432[40] = |(datain[151:148] ^ 14);
  assign w432[41] = |(datain[147:144] ^ 8);
  assign w432[42] = |(datain[143:140] ^ 4);
  assign w432[43] = |(datain[139:136] ^ 8);
  assign w432[44] = |(datain[135:132] ^ 0);
  assign w432[45] = |(datain[131:128] ^ 0);
  assign w432[46] = |(datain[127:124] ^ 7);
  assign w432[47] = |(datain[123:120] ^ 2);
  assign w432[48] = |(datain[119:116] ^ 1);
  assign w432[49] = |(datain[115:112] ^ 10);
  assign w432[50] = |(datain[111:108] ^ 11);
  assign w432[51] = |(datain[107:104] ^ 9);
  assign w432[52] = |(datain[103:100] ^ 0);
  assign w432[53] = |(datain[99:96] ^ 3);
  assign w432[54] = |(datain[95:92] ^ 0);
  assign w432[55] = |(datain[91:88] ^ 0);
  assign w432[56] = |(datain[87:84] ^ 11);
  assign w432[57] = |(datain[83:80] ^ 10);
  assign w432[58] = |(datain[79:76] ^ 8);
  assign w432[59] = |(datain[75:72] ^ 6);
  assign w432[60] = |(datain[71:68] ^ 0);
  assign w432[61] = |(datain[67:64] ^ 5);
  assign w432[62] = |(datain[63:60] ^ 11);
  assign w432[63] = |(datain[59:56] ^ 4);
  assign w432[64] = |(datain[55:52] ^ 4);
  assign w432[65] = |(datain[51:48] ^ 0);
  assign w432[66] = |(datain[47:44] ^ 14);
  assign w432[67] = |(datain[43:40] ^ 8);
  assign w432[68] = |(datain[39:36] ^ 3);
  assign w432[69] = |(datain[35:32] ^ 11);
  assign w432[70] = |(datain[31:28] ^ 0);
  assign w432[71] = |(datain[27:24] ^ 0);
  assign w432[72] = |(datain[23:20] ^ 7);
  assign w432[73] = |(datain[19:16] ^ 2);
  assign comp[432] = ~(|w432);
  wire [34-1:0] w433;
  assign w433[0] = |(datain[311:308] ^ 0);
  assign w433[1] = |(datain[307:304] ^ 1);
  assign w433[2] = |(datain[303:300] ^ 0);
  assign w433[3] = |(datain[299:296] ^ 1);
  assign w433[4] = |(datain[295:292] ^ 8);
  assign w433[5] = |(datain[291:288] ^ 13);
  assign w433[6] = |(datain[287:284] ^ 11);
  assign w433[7] = |(datain[283:280] ^ 14);
  assign w433[8] = |(datain[279:276] ^ 1);
  assign w433[9] = |(datain[275:272] ^ 5);
  assign w433[10] = |(datain[271:268] ^ 0);
  assign w433[11] = |(datain[267:264] ^ 1);
  assign w433[12] = |(datain[263:260] ^ 11);
  assign w433[13] = |(datain[259:256] ^ 9);
  assign w433[14] = |(datain[255:252] ^ 12);
  assign w433[15] = |(datain[251:248] ^ 3);
  assign w433[16] = |(datain[247:244] ^ 0);
  assign w433[17] = |(datain[243:240] ^ 1);
  assign w433[18] = |(datain[239:236] ^ 10);
  assign w433[19] = |(datain[235:232] ^ 13);
  assign w433[20] = |(datain[231:228] ^ 8);
  assign w433[21] = |(datain[227:224] ^ 11);
  assign w433[22] = |(datain[223:220] ^ 13);
  assign w433[23] = |(datain[219:216] ^ 0);
  assign w433[24] = |(datain[215:212] ^ 3);
  assign w433[25] = |(datain[211:208] ^ 1);
  assign w433[26] = |(datain[207:204] ^ 1);
  assign w433[27] = |(datain[203:200] ^ 5);
  assign w433[28] = |(datain[199:196] ^ 4);
  assign w433[29] = |(datain[195:192] ^ 7);
  assign w433[30] = |(datain[191:188] ^ 14);
  assign w433[31] = |(datain[187:184] ^ 2);
  assign w433[32] = |(datain[183:180] ^ 15);
  assign w433[33] = |(datain[179:176] ^ 11);
  assign comp[433] = ~(|w433);
  wire [40-1:0] w434;
  assign w434[0] = |(datain[311:308] ^ 11);
  assign w434[1] = |(datain[307:304] ^ 4);
  assign w434[2] = |(datain[303:300] ^ 4);
  assign w434[3] = |(datain[299:296] ^ 0);
  assign w434[4] = |(datain[295:292] ^ 8);
  assign w434[5] = |(datain[291:288] ^ 11);
  assign w434[6] = |(datain[287:284] ^ 9);
  assign w434[7] = |(datain[283:280] ^ 12);
  assign w434[8] = |(datain[279:276] ^ 3);
  assign w434[9] = |(datain[275:272] ^ 5);
  assign w434[10] = |(datain[271:268] ^ 0);
  assign w434[11] = |(datain[267:264] ^ 4);
  assign w434[12] = |(datain[263:260] ^ 11);
  assign w434[13] = |(datain[259:256] ^ 9);
  assign w434[14] = |(datain[255:252] ^ 14);
  assign w434[15] = |(datain[251:248] ^ 6);
  assign w434[16] = |(datain[247:244] ^ 0);
  assign w434[17] = |(datain[243:240] ^ 2);
  assign w434[18] = |(datain[239:236] ^ 8);
  assign w434[19] = |(datain[235:232] ^ 13);
  assign w434[20] = |(datain[231:228] ^ 9);
  assign w434[21] = |(datain[227:224] ^ 4);
  assign w434[22] = |(datain[223:220] ^ 0);
  assign w434[23] = |(datain[219:216] ^ 14);
  assign w434[24] = |(datain[215:212] ^ 0);
  assign w434[25] = |(datain[211:208] ^ 1);
  assign w434[26] = |(datain[207:204] ^ 12);
  assign w434[27] = |(datain[203:200] ^ 13);
  assign w434[28] = |(datain[199:196] ^ 2);
  assign w434[29] = |(datain[195:192] ^ 1);
  assign w434[30] = |(datain[191:188] ^ 14);
  assign w434[31] = |(datain[187:184] ^ 8);
  assign w434[32] = |(datain[183:180] ^ 13);
  assign w434[33] = |(datain[179:176] ^ 6);
  assign w434[34] = |(datain[175:172] ^ 15);
  assign w434[35] = |(datain[171:168] ^ 15);
  assign w434[36] = |(datain[167:164] ^ 14);
  assign w434[37] = |(datain[163:160] ^ 8);
  assign w434[38] = |(datain[159:156] ^ 11);
  assign w434[39] = |(datain[155:152] ^ 14);
  assign comp[434] = ~(|w434);
  wire [44-1:0] w435;
  assign w435[0] = |(datain[311:308] ^ 8);
  assign w435[1] = |(datain[307:304] ^ 13);
  assign w435[2] = |(datain[303:300] ^ 11);
  assign w435[3] = |(datain[299:296] ^ 6);
  assign w435[4] = |(datain[295:292] ^ 2);
  assign w435[5] = |(datain[291:288] ^ 7);
  assign w435[6] = |(datain[287:284] ^ 0);
  assign w435[7] = |(datain[283:280] ^ 1);
  assign w435[8] = |(datain[279:276] ^ 5);
  assign w435[9] = |(datain[275:272] ^ 6);
  assign w435[10] = |(datain[271:268] ^ 8);
  assign w435[11] = |(datain[267:264] ^ 11);
  assign w435[12] = |(datain[263:260] ^ 9);
  assign w435[13] = |(datain[259:256] ^ 6);
  assign w435[14] = |(datain[255:252] ^ 15);
  assign w435[15] = |(datain[251:248] ^ 2);
  assign w435[16] = |(datain[247:244] ^ 0);
  assign w435[17] = |(datain[243:240] ^ 1);
  assign w435[18] = |(datain[239:236] ^ 11);
  assign w435[19] = |(datain[235:232] ^ 9);
  assign w435[20] = |(datain[231:228] ^ 6);
  assign w435[21] = |(datain[227:224] ^ 0);
  assign w435[22] = |(datain[223:220] ^ 0);
  assign w435[23] = |(datain[219:216] ^ 0);
  assign w435[24] = |(datain[215:212] ^ 8);
  assign w435[25] = |(datain[211:208] ^ 11);
  assign w435[26] = |(datain[207:204] ^ 15);
  assign w435[27] = |(datain[203:200] ^ 14);
  assign w435[28] = |(datain[199:196] ^ 15);
  assign w435[29] = |(datain[195:192] ^ 12);
  assign w435[30] = |(datain[191:188] ^ 10);
  assign w435[31] = |(datain[187:184] ^ 13);
  assign w435[32] = |(datain[183:180] ^ 3);
  assign w435[33] = |(datain[179:176] ^ 3);
  assign w435[34] = |(datain[175:172] ^ 12);
  assign w435[35] = |(datain[171:168] ^ 2);
  assign w435[36] = |(datain[167:164] ^ 10);
  assign w435[37] = |(datain[163:160] ^ 11);
  assign w435[38] = |(datain[159:156] ^ 14);
  assign w435[39] = |(datain[155:152] ^ 2);
  assign w435[40] = |(datain[151:148] ^ 15);
  assign w435[41] = |(datain[147:144] ^ 10);
  assign w435[42] = |(datain[143:140] ^ 12);
  assign w435[43] = |(datain[139:136] ^ 3);
  assign comp[435] = ~(|w435);
  wire [44-1:0] w436;
  assign w436[0] = |(datain[311:308] ^ 8);
  assign w436[1] = |(datain[307:304] ^ 13);
  assign w436[2] = |(datain[303:300] ^ 11);
  assign w436[3] = |(datain[299:296] ^ 6);
  assign w436[4] = |(datain[295:292] ^ 3);
  assign w436[5] = |(datain[291:288] ^ 13);
  assign w436[6] = |(datain[287:284] ^ 0);
  assign w436[7] = |(datain[283:280] ^ 1);
  assign w436[8] = |(datain[279:276] ^ 5);
  assign w436[9] = |(datain[275:272] ^ 6);
  assign w436[10] = |(datain[271:268] ^ 8);
  assign w436[11] = |(datain[267:264] ^ 11);
  assign w436[12] = |(datain[263:260] ^ 9);
  assign w436[13] = |(datain[259:256] ^ 6);
  assign w436[14] = |(datain[255:252] ^ 1);
  assign w436[15] = |(datain[251:248] ^ 8);
  assign w436[16] = |(datain[247:244] ^ 0);
  assign w436[17] = |(datain[243:240] ^ 2);
  assign w436[18] = |(datain[239:236] ^ 11);
  assign w436[19] = |(datain[235:232] ^ 9);
  assign w436[20] = |(datain[231:228] ^ 6);
  assign w436[21] = |(datain[227:224] ^ 13);
  assign w436[22] = |(datain[223:220] ^ 0);
  assign w436[23] = |(datain[219:216] ^ 0);
  assign w436[24] = |(datain[215:212] ^ 8);
  assign w436[25] = |(datain[211:208] ^ 11);
  assign w436[26] = |(datain[207:204] ^ 15);
  assign w436[27] = |(datain[203:200] ^ 14);
  assign w436[28] = |(datain[199:196] ^ 15);
  assign w436[29] = |(datain[195:192] ^ 12);
  assign w436[30] = |(datain[191:188] ^ 10);
  assign w436[31] = |(datain[187:184] ^ 13);
  assign w436[32] = |(datain[183:180] ^ 3);
  assign w436[33] = |(datain[179:176] ^ 3);
  assign w436[34] = |(datain[175:172] ^ 12);
  assign w436[35] = |(datain[171:168] ^ 2);
  assign w436[36] = |(datain[167:164] ^ 10);
  assign w436[37] = |(datain[163:160] ^ 11);
  assign w436[38] = |(datain[159:156] ^ 14);
  assign w436[39] = |(datain[155:152] ^ 2);
  assign w436[40] = |(datain[151:148] ^ 15);
  assign w436[41] = |(datain[147:144] ^ 10);
  assign w436[42] = |(datain[143:140] ^ 12);
  assign w436[43] = |(datain[139:136] ^ 3);
  assign comp[436] = ~(|w436);
  wire [48-1:0] w437;
  assign w437[0] = |(datain[311:308] ^ 6);
  assign w437[1] = |(datain[307:304] ^ 0);
  assign w437[2] = |(datain[303:300] ^ 14);
  assign w437[3] = |(datain[299:296] ^ 8);
  assign w437[4] = |(datain[295:292] ^ 0);
  assign w437[5] = |(datain[291:288] ^ 0);
  assign w437[6] = |(datain[287:284] ^ 0);
  assign w437[7] = |(datain[283:280] ^ 0);
  assign w437[8] = |(datain[279:276] ^ 5);
  assign w437[9] = |(datain[275:272] ^ 8);
  assign w437[10] = |(datain[271:268] ^ 2);
  assign w437[11] = |(datain[267:264] ^ 13);
  assign w437[12] = |(datain[263:260] ^ 8);
  assign w437[13] = |(datain[259:256] ^ 11);
  assign w437[14] = |(datain[255:252] ^ 0);
  assign w437[15] = |(datain[251:248] ^ 1);
  assign w437[16] = |(datain[247:244] ^ 9);
  assign w437[17] = |(datain[243:240] ^ 5);
  assign w437[18] = |(datain[239:236] ^ 8);
  assign w437[19] = |(datain[235:232] ^ 13);
  assign w437[20] = |(datain[231:228] ^ 11);
  assign w437[21] = |(datain[227:224] ^ 6);
  assign w437[22] = |(datain[223:220] ^ 10);
  assign w437[23] = |(datain[219:216] ^ 12);
  assign w437[24] = |(datain[215:212] ^ 0);
  assign w437[25] = |(datain[211:208] ^ 1);
  assign w437[26] = |(datain[207:204] ^ 14);
  assign w437[27] = |(datain[203:200] ^ 8);
  assign w437[28] = |(datain[199:196] ^ 0);
  assign w437[29] = |(datain[195:192] ^ 2);
  assign w437[30] = |(datain[191:188] ^ 0);
  assign w437[31] = |(datain[187:184] ^ 0);
  assign w437[32] = |(datain[183:180] ^ 14);
  assign w437[33] = |(datain[179:176] ^ 11);
  assign w437[34] = |(datain[175:172] ^ 1);
  assign w437[35] = |(datain[171:168] ^ 3);
  assign w437[36] = |(datain[167:164] ^ 11);
  assign w437[37] = |(datain[163:160] ^ 9);
  assign w437[38] = |(datain[159:156] ^ 1);
  assign w437[39] = |(datain[155:152] ^ 7);
  assign w437[40] = |(datain[151:148] ^ 0);
  assign w437[41] = |(datain[147:144] ^ 1);
  assign w437[42] = |(datain[143:140] ^ 8);
  assign w437[43] = |(datain[139:136] ^ 11);
  assign w437[44] = |(datain[135:132] ^ 15);
  assign w437[45] = |(datain[131:128] ^ 14);
  assign w437[46] = |(datain[127:124] ^ 11);
  assign w437[47] = |(datain[123:120] ^ 10);
  assign comp[437] = ~(|w437);
  wire [46-1:0] w438;
  assign w438[0] = |(datain[311:308] ^ 14);
  assign w438[1] = |(datain[307:304] ^ 8);
  assign w438[2] = |(datain[303:300] ^ 0);
  assign w438[3] = |(datain[299:296] ^ 0);
  assign w438[4] = |(datain[295:292] ^ 0);
  assign w438[5] = |(datain[291:288] ^ 0);
  assign w438[6] = |(datain[287:284] ^ 5);
  assign w438[7] = |(datain[283:280] ^ 11);
  assign w438[8] = |(datain[279:276] ^ 8);
  assign w438[9] = |(datain[275:272] ^ 1);
  assign w438[10] = |(datain[271:268] ^ 14);
  assign w438[11] = |(datain[267:264] ^ 11);
  assign w438[12] = |(datain[263:260] ^ 0);
  assign w438[13] = |(datain[259:256] ^ 10);
  assign w438[14] = |(datain[255:252] ^ 0);
  assign w438[15] = |(datain[251:248] ^ 1);
  assign w438[16] = |(datain[247:244] ^ 8);
  assign w438[17] = |(datain[243:240] ^ 13);
  assign w438[18] = |(datain[239:236] ^ 11);
  assign w438[19] = |(datain[235:232] ^ 7);
  assign w438[20] = |(datain[231:228] ^ 2);
  assign w438[21] = |(datain[227:224] ^ 11);
  assign w438[22] = |(datain[223:220] ^ 0);
  assign w438[23] = |(datain[219:216] ^ 1);
  assign w438[24] = |(datain[215:212] ^ 14);
  assign w438[25] = |(datain[211:208] ^ 8);
  assign w438[26] = |(datain[207:204] ^ 0);
  assign w438[27] = |(datain[203:200] ^ 2);
  assign w438[28] = |(datain[199:196] ^ 0);
  assign w438[29] = |(datain[195:192] ^ 0);
  assign w438[30] = |(datain[191:188] ^ 14);
  assign w438[31] = |(datain[187:184] ^ 11);
  assign w438[32] = |(datain[183:180] ^ 1);
  assign w438[33] = |(datain[179:176] ^ 3);
  assign w438[34] = |(datain[175:172] ^ 11);
  assign w438[35] = |(datain[171:168] ^ 9);
  assign w438[36] = |(datain[167:164] ^ 1);
  assign w438[37] = |(datain[163:160] ^ 8);
  assign w438[38] = |(datain[159:156] ^ 0);
  assign w438[39] = |(datain[155:152] ^ 1);
  assign w438[40] = |(datain[151:148] ^ 8);
  assign w438[41] = |(datain[147:144] ^ 11);
  assign w438[42] = |(datain[143:140] ^ 15);
  assign w438[43] = |(datain[139:136] ^ 14);
  assign w438[44] = |(datain[135:132] ^ 11);
  assign w438[45] = |(datain[131:128] ^ 10);
  assign comp[438] = ~(|w438);
  wire [46-1:0] w439;
  assign w439[0] = |(datain[311:308] ^ 14);
  assign w439[1] = |(datain[307:304] ^ 8);
  assign w439[2] = |(datain[303:300] ^ 0);
  assign w439[3] = |(datain[299:296] ^ 0);
  assign w439[4] = |(datain[295:292] ^ 0);
  assign w439[5] = |(datain[291:288] ^ 0);
  assign w439[6] = |(datain[287:284] ^ 5);
  assign w439[7] = |(datain[283:280] ^ 8);
  assign w439[8] = |(datain[279:276] ^ 2);
  assign w439[9] = |(datain[275:272] ^ 13);
  assign w439[10] = |(datain[271:268] ^ 0);
  assign w439[11] = |(datain[267:264] ^ 10);
  assign w439[12] = |(datain[263:260] ^ 0);
  assign w439[13] = |(datain[259:256] ^ 1);
  assign w439[14] = |(datain[255:252] ^ 9);
  assign w439[15] = |(datain[251:248] ^ 5);
  assign w439[16] = |(datain[247:244] ^ 8);
  assign w439[17] = |(datain[243:240] ^ 13);
  assign w439[18] = |(datain[239:236] ^ 11);
  assign w439[19] = |(datain[235:232] ^ 6);
  assign w439[20] = |(datain[231:228] ^ 2);
  assign w439[21] = |(datain[227:224] ^ 11);
  assign w439[22] = |(datain[223:220] ^ 0);
  assign w439[23] = |(datain[219:216] ^ 1);
  assign w439[24] = |(datain[215:212] ^ 14);
  assign w439[25] = |(datain[211:208] ^ 8);
  assign w439[26] = |(datain[207:204] ^ 0);
  assign w439[27] = |(datain[203:200] ^ 2);
  assign w439[28] = |(datain[199:196] ^ 0);
  assign w439[29] = |(datain[195:192] ^ 0);
  assign w439[30] = |(datain[191:188] ^ 14);
  assign w439[31] = |(datain[187:184] ^ 11);
  assign w439[32] = |(datain[183:180] ^ 1);
  assign w439[33] = |(datain[179:176] ^ 3);
  assign w439[34] = |(datain[175:172] ^ 11);
  assign w439[35] = |(datain[171:168] ^ 9);
  assign w439[36] = |(datain[167:164] ^ 1);
  assign w439[37] = |(datain[163:160] ^ 12);
  assign w439[38] = |(datain[159:156] ^ 0);
  assign w439[39] = |(datain[155:152] ^ 1);
  assign w439[40] = |(datain[151:148] ^ 8);
  assign w439[41] = |(datain[147:144] ^ 11);
  assign w439[42] = |(datain[143:140] ^ 15);
  assign w439[43] = |(datain[139:136] ^ 14);
  assign w439[44] = |(datain[135:132] ^ 11);
  assign w439[45] = |(datain[131:128] ^ 10);
  assign comp[439] = ~(|w439);
  wire [48-1:0] w440;
  assign w440[0] = |(datain[311:308] ^ 6);
  assign w440[1] = |(datain[307:304] ^ 0);
  assign w440[2] = |(datain[303:300] ^ 14);
  assign w440[3] = |(datain[299:296] ^ 8);
  assign w440[4] = |(datain[295:292] ^ 0);
  assign w440[5] = |(datain[291:288] ^ 0);
  assign w440[6] = |(datain[287:284] ^ 0);
  assign w440[7] = |(datain[283:280] ^ 0);
  assign w440[8] = |(datain[279:276] ^ 5);
  assign w440[9] = |(datain[275:272] ^ 8);
  assign w440[10] = |(datain[271:268] ^ 2);
  assign w440[11] = |(datain[267:264] ^ 13);
  assign w440[12] = |(datain[263:260] ^ 0);
  assign w440[13] = |(datain[259:256] ^ 10);
  assign w440[14] = |(datain[255:252] ^ 0);
  assign w440[15] = |(datain[251:248] ^ 1);
  assign w440[16] = |(datain[247:244] ^ 9);
  assign w440[17] = |(datain[243:240] ^ 5);
  assign w440[18] = |(datain[239:236] ^ 8);
  assign w440[19] = |(datain[235:232] ^ 13);
  assign w440[20] = |(datain[231:228] ^ 11);
  assign w440[21] = |(datain[227:224] ^ 6);
  assign w440[22] = |(datain[223:220] ^ 2);
  assign w440[23] = |(datain[219:216] ^ 11);
  assign w440[24] = |(datain[215:212] ^ 0);
  assign w440[25] = |(datain[211:208] ^ 1);
  assign w440[26] = |(datain[207:204] ^ 14);
  assign w440[27] = |(datain[203:200] ^ 8);
  assign w440[28] = |(datain[199:196] ^ 0);
  assign w440[29] = |(datain[195:192] ^ 2);
  assign w440[30] = |(datain[191:188] ^ 0);
  assign w440[31] = |(datain[187:184] ^ 0);
  assign w440[32] = |(datain[183:180] ^ 14);
  assign w440[33] = |(datain[179:176] ^ 11);
  assign w440[34] = |(datain[175:172] ^ 1);
  assign w440[35] = |(datain[171:168] ^ 3);
  assign w440[36] = |(datain[167:164] ^ 11);
  assign w440[37] = |(datain[163:160] ^ 9);
  assign w440[38] = |(datain[159:156] ^ 1);
  assign w440[39] = |(datain[155:152] ^ 14);
  assign w440[40] = |(datain[151:148] ^ 0);
  assign w440[41] = |(datain[147:144] ^ 1);
  assign w440[42] = |(datain[143:140] ^ 8);
  assign w440[43] = |(datain[139:136] ^ 11);
  assign w440[44] = |(datain[135:132] ^ 15);
  assign w440[45] = |(datain[131:128] ^ 14);
  assign w440[46] = |(datain[127:124] ^ 11);
  assign w440[47] = |(datain[123:120] ^ 10);
  assign comp[440] = ~(|w440);
  wire [76-1:0] w441;
  assign w441[0] = |(datain[311:308] ^ 0);
  assign w441[1] = |(datain[307:304] ^ 2);
  assign w441[2] = |(datain[303:300] ^ 10);
  assign w441[3] = |(datain[299:296] ^ 3);
  assign w441[4] = |(datain[295:292] ^ 0);
  assign w441[5] = |(datain[291:288] ^ 5);
  assign w441[6] = |(datain[287:284] ^ 0);
  assign w441[7] = |(datain[283:280] ^ 0);
  assign w441[8] = |(datain[279:276] ^ 1);
  assign w441[9] = |(datain[275:272] ^ 14);
  assign w441[10] = |(datain[271:268] ^ 8);
  assign w441[11] = |(datain[267:264] ^ 11);
  assign w441[12] = |(datain[263:260] ^ 1);
  assign w441[13] = |(datain[259:256] ^ 6);
  assign w441[14] = |(datain[255:252] ^ 8);
  assign w441[15] = |(datain[251:248] ^ 2);
  assign w441[16] = |(datain[247:244] ^ 0);
  assign w441[17] = |(datain[243:240] ^ 2);
  assign w441[18] = |(datain[239:236] ^ 8);
  assign w441[19] = |(datain[235:232] ^ 3);
  assign w441[20] = |(datain[231:228] ^ 14);
  assign w441[21] = |(datain[227:224] ^ 2);
  assign w441[22] = |(datain[223:220] ^ 0);
  assign w441[23] = |(datain[219:216] ^ 15);
  assign w441[24] = |(datain[215:212] ^ 11);
  assign w441[25] = |(datain[211:208] ^ 9);
  assign w441[26] = |(datain[207:204] ^ 9);
  assign w441[27] = |(datain[203:200] ^ 0);
  assign w441[28] = |(datain[199:196] ^ 0);
  assign w441[29] = |(datain[195:192] ^ 2);
  assign w441[30] = |(datain[191:188] ^ 8);
  assign w441[31] = |(datain[187:184] ^ 12);
  assign w441[32] = |(datain[183:180] ^ 13);
  assign w441[33] = |(datain[179:176] ^ 8);
  assign w441[34] = |(datain[175:172] ^ 4);
  assign w441[35] = |(datain[171:168] ^ 8);
  assign w441[36] = |(datain[167:164] ^ 8);
  assign w441[37] = |(datain[163:160] ^ 14);
  assign w441[38] = |(datain[159:156] ^ 13);
  assign w441[39] = |(datain[155:152] ^ 8);
  assign w441[40] = |(datain[151:148] ^ 11);
  assign w441[41] = |(datain[147:144] ^ 4);
  assign w441[42] = |(datain[143:140] ^ 4);
  assign w441[43] = |(datain[139:136] ^ 0);
  assign w441[44] = |(datain[135:132] ^ 14);
  assign w441[45] = |(datain[131:128] ^ 8);
  assign w441[46] = |(datain[127:124] ^ 10);
  assign w441[47] = |(datain[123:120] ^ 14);
  assign w441[48] = |(datain[119:116] ^ 0);
  assign w441[49] = |(datain[115:112] ^ 0);
  assign w441[50] = |(datain[111:108] ^ 1);
  assign w441[51] = |(datain[107:104] ^ 15);
  assign w441[52] = |(datain[103:100] ^ 7);
  assign w441[53] = |(datain[99:96] ^ 2);
  assign w441[54] = |(datain[95:92] ^ 5);
  assign w441[55] = |(datain[91:88] ^ 7);
  assign w441[56] = |(datain[87:84] ^ 3);
  assign w441[57] = |(datain[83:80] ^ 3);
  assign w441[58] = |(datain[79:76] ^ 13);
  assign w441[59] = |(datain[75:72] ^ 2);
  assign w441[60] = |(datain[71:68] ^ 10);
  assign w441[61] = |(datain[67:64] ^ 1);
  assign w441[62] = |(datain[63:60] ^ 8);
  assign w441[63] = |(datain[59:56] ^ 4);
  assign w441[64] = |(datain[55:52] ^ 0);
  assign w441[65] = |(datain[51:48] ^ 2);
  assign w441[66] = |(datain[47:44] ^ 4);
  assign w441[67] = |(datain[43:40] ^ 8);
  assign w441[68] = |(datain[39:36] ^ 11);
  assign w441[69] = |(datain[35:32] ^ 9);
  assign w441[70] = |(datain[31:28] ^ 2);
  assign w441[71] = |(datain[27:24] ^ 0);
  assign w441[72] = |(datain[23:20] ^ 0);
  assign w441[73] = |(datain[19:16] ^ 0);
  assign w441[74] = |(datain[15:12] ^ 15);
  assign w441[75] = |(datain[11:8] ^ 7);
  assign comp[441] = ~(|w441);
  wire [42-1:0] w442;
  assign w442[0] = |(datain[311:308] ^ 11);
  assign w442[1] = |(datain[307:304] ^ 4);
  assign w442[2] = |(datain[303:300] ^ 3);
  assign w442[3] = |(datain[299:296] ^ 15);
  assign w442[4] = |(datain[295:292] ^ 11);
  assign w442[5] = |(datain[291:288] ^ 9);
  assign w442[6] = |(datain[287:284] ^ 1);
  assign w442[7] = |(datain[283:280] ^ 5);
  assign w442[8] = |(datain[279:276] ^ 0);
  assign w442[9] = |(datain[275:272] ^ 1);
  assign w442[10] = |(datain[271:268] ^ 8);
  assign w442[11] = |(datain[267:264] ^ 13);
  assign w442[12] = |(datain[263:260] ^ 9);
  assign w442[13] = |(datain[259:256] ^ 6);
  assign w442[14] = |(datain[255:252] ^ 0);
  assign w442[15] = |(datain[251:248] ^ 3);
  assign w442[16] = |(datain[247:244] ^ 0);
  assign w442[17] = |(datain[243:240] ^ 1);
  assign w442[18] = |(datain[239:236] ^ 15);
  assign w442[19] = |(datain[235:232] ^ 14);
  assign w442[20] = |(datain[231:228] ^ 12);
  assign w442[21] = |(datain[227:224] ^ 4);
  assign w442[22] = |(datain[223:220] ^ 12);
  assign w442[23] = |(datain[219:216] ^ 13);
  assign w442[24] = |(datain[215:212] ^ 2);
  assign w442[25] = |(datain[211:208] ^ 1);
  assign w442[26] = |(datain[207:204] ^ 11);
  assign w442[27] = |(datain[203:200] ^ 8);
  assign w442[28] = |(datain[199:196] ^ 0);
  assign w442[29] = |(datain[195:192] ^ 1);
  assign w442[30] = |(datain[191:188] ^ 5);
  assign w442[31] = |(datain[187:184] ^ 7);
  assign w442[32] = |(datain[183:180] ^ 3);
  assign w442[33] = |(datain[179:176] ^ 14);
  assign w442[34] = |(datain[175:172] ^ 8);
  assign w442[35] = |(datain[171:168] ^ 11);
  assign w442[36] = |(datain[167:164] ^ 8);
  assign w442[37] = |(datain[163:160] ^ 14);
  assign w442[38] = |(datain[159:156] ^ 3);
  assign w442[39] = |(datain[155:152] ^ 1);
  assign w442[40] = |(datain[151:148] ^ 0);
  assign w442[41] = |(datain[147:144] ^ 2);
  assign comp[442] = ~(|w442);
  wire [76-1:0] w443;
  assign w443[0] = |(datain[311:308] ^ 8);
  assign w443[1] = |(datain[307:304] ^ 6);
  assign w443[2] = |(datain[303:300] ^ 6);
  assign w443[3] = |(datain[299:296] ^ 1);
  assign w443[4] = |(datain[295:292] ^ 0);
  assign w443[5] = |(datain[291:288] ^ 4);
  assign w443[6] = |(datain[287:284] ^ 8);
  assign w443[7] = |(datain[283:280] ^ 13);
  assign w443[8] = |(datain[279:276] ^ 9);
  assign w443[9] = |(datain[275:272] ^ 6);
  assign w443[10] = |(datain[271:268] ^ 0);
  assign w443[11] = |(datain[267:264] ^ 2);
  assign w443[12] = |(datain[263:260] ^ 0);
  assign w443[13] = |(datain[259:256] ^ 3);
  assign w443[14] = |(datain[255:252] ^ 11);
  assign w443[15] = |(datain[251:248] ^ 4);
  assign w443[16] = |(datain[247:244] ^ 4);
  assign w443[17] = |(datain[243:240] ^ 0);
  assign w443[18] = |(datain[239:236] ^ 11);
  assign w443[19] = |(datain[235:232] ^ 9);
  assign w443[20] = |(datain[231:228] ^ 6);
  assign w443[21] = |(datain[227:224] ^ 15);
  assign w443[22] = |(datain[223:220] ^ 0);
  assign w443[23] = |(datain[219:216] ^ 1);
  assign w443[24] = |(datain[215:212] ^ 12);
  assign w443[25] = |(datain[211:208] ^ 13);
  assign w443[26] = |(datain[207:204] ^ 2);
  assign w443[27] = |(datain[203:200] ^ 1);
  assign w443[28] = |(datain[199:196] ^ 11);
  assign w443[29] = |(datain[195:192] ^ 8);
  assign w443[30] = |(datain[191:188] ^ 0);
  assign w443[31] = |(datain[187:184] ^ 0);
  assign w443[32] = |(datain[183:180] ^ 4);
  assign w443[33] = |(datain[179:176] ^ 2);
  assign w443[34] = |(datain[175:172] ^ 2);
  assign w443[35] = |(datain[171:168] ^ 11);
  assign w443[36] = |(datain[167:164] ^ 13);
  assign w443[37] = |(datain[163:160] ^ 2);
  assign w443[38] = |(datain[159:156] ^ 2);
  assign w443[39] = |(datain[155:152] ^ 11);
  assign w443[40] = |(datain[151:148] ^ 12);
  assign w443[41] = |(datain[147:144] ^ 9);
  assign w443[42] = |(datain[143:140] ^ 12);
  assign w443[43] = |(datain[139:136] ^ 13);
  assign w443[44] = |(datain[135:132] ^ 2);
  assign w443[45] = |(datain[131:128] ^ 1);
  assign w443[46] = |(datain[127:124] ^ 8);
  assign w443[47] = |(datain[123:120] ^ 13);
  assign w443[48] = |(datain[119:116] ^ 9);
  assign w443[49] = |(datain[115:112] ^ 6);
  assign w443[50] = |(datain[111:108] ^ 6);
  assign w443[51] = |(datain[107:104] ^ 0);
  assign w443[52] = |(datain[103:100] ^ 0);
  assign w443[53] = |(datain[99:96] ^ 4);
  assign w443[54] = |(datain[95:92] ^ 11);
  assign w443[55] = |(datain[91:88] ^ 4);
  assign w443[56] = |(datain[87:84] ^ 4);
  assign w443[57] = |(datain[83:80] ^ 0);
  assign w443[58] = |(datain[79:76] ^ 11);
  assign w443[59] = |(datain[75:72] ^ 9);
  assign w443[60] = |(datain[71:68] ^ 0);
  assign w443[61] = |(datain[67:64] ^ 3);
  assign w443[62] = |(datain[63:60] ^ 0);
  assign w443[63] = |(datain[59:56] ^ 0);
  assign w443[64] = |(datain[55:52] ^ 12);
  assign w443[65] = |(datain[51:48] ^ 13);
  assign w443[66] = |(datain[47:44] ^ 2);
  assign w443[67] = |(datain[43:40] ^ 1);
  assign w443[68] = |(datain[39:36] ^ 14);
  assign w443[69] = |(datain[35:32] ^ 8);
  assign w443[70] = |(datain[31:28] ^ 4);
  assign w443[71] = |(datain[27:24] ^ 0);
  assign w443[72] = |(datain[23:20] ^ 0);
  assign w443[73] = |(datain[19:16] ^ 0);
  assign w443[74] = |(datain[15:12] ^ 5);
  assign w443[75] = |(datain[11:8] ^ 10);
  assign comp[443] = ~(|w443);
  wire [28-1:0] w444;
  assign w444[0] = |(datain[311:308] ^ 8);
  assign w444[1] = |(datain[307:304] ^ 3);
  assign w444[2] = |(datain[303:300] ^ 2);
  assign w444[3] = |(datain[299:296] ^ 14);
  assign w444[4] = |(datain[295:292] ^ 1);
  assign w444[5] = |(datain[291:288] ^ 3);
  assign w444[6] = |(datain[287:284] ^ 0);
  assign w444[7] = |(datain[283:280] ^ 4);
  assign w444[8] = |(datain[279:276] ^ 0);
  assign w444[9] = |(datain[275:272] ^ 2);
  assign w444[10] = |(datain[271:268] ^ 12);
  assign w444[11] = |(datain[267:264] ^ 13);
  assign w444[12] = |(datain[263:260] ^ 1);
  assign w444[13] = |(datain[259:256] ^ 2);
  assign w444[14] = |(datain[255:252] ^ 11);
  assign w444[15] = |(datain[251:248] ^ 1);
  assign w444[16] = |(datain[247:244] ^ 0);
  assign w444[17] = |(datain[243:240] ^ 6);
  assign w444[18] = |(datain[239:236] ^ 13);
  assign w444[19] = |(datain[235:232] ^ 3);
  assign w444[20] = |(datain[231:228] ^ 14);
  assign w444[21] = |(datain[227:224] ^ 0);
  assign w444[22] = |(datain[223:220] ^ 8);
  assign w444[23] = |(datain[219:216] ^ 14);
  assign w444[24] = |(datain[215:212] ^ 12);
  assign w444[25] = |(datain[211:208] ^ 0);
  assign w444[26] = |(datain[207:204] ^ 11);
  assign w444[27] = |(datain[203:200] ^ 15);
  assign comp[444] = ~(|w444);
  wire [32-1:0] w445;
  assign w445[0] = |(datain[311:308] ^ 1);
  assign w445[1] = |(datain[307:304] ^ 3);
  assign w445[2] = |(datain[303:300] ^ 5);
  assign w445[3] = |(datain[299:296] ^ 8);
  assign w445[4] = |(datain[295:292] ^ 11);
  assign w445[5] = |(datain[291:288] ^ 1);
  assign w445[6] = |(datain[287:284] ^ 0);
  assign w445[7] = |(datain[283:280] ^ 1);
  assign w445[8] = |(datain[279:276] ^ 11);
  assign w445[9] = |(datain[275:272] ^ 11);
  assign w445[10] = |(datain[271:268] ^ 0);
  assign w445[11] = |(datain[267:264] ^ 0);
  assign w445[12] = |(datain[263:260] ^ 0);
  assign w445[13] = |(datain[259:256] ^ 4);
  assign w445[14] = |(datain[255:252] ^ 12);
  assign w445[15] = |(datain[251:248] ^ 13);
  assign w445[16] = |(datain[247:244] ^ 1);
  assign w445[17] = |(datain[243:240] ^ 3);
  assign w445[18] = |(datain[239:236] ^ 0);
  assign w445[19] = |(datain[235:232] ^ 14);
  assign w445[20] = |(datain[231:228] ^ 1);
  assign w445[21] = |(datain[227:224] ^ 15);
  assign w445[22] = |(datain[223:220] ^ 11);
  assign w445[23] = |(datain[219:216] ^ 14);
  assign w445[24] = |(datain[215:212] ^ 9);
  assign w445[25] = |(datain[211:208] ^ 11);
  assign w445[26] = |(datain[207:204] ^ 0);
  assign w445[27] = |(datain[203:200] ^ 3);
  assign w445[28] = |(datain[199:196] ^ 8);
  assign w445[29] = |(datain[195:192] ^ 11);
  assign w445[30] = |(datain[191:188] ^ 15);
  assign w445[31] = |(datain[187:184] ^ 11);
  assign comp[445] = ~(|w445);
  wire [30-1:0] w446;
  assign w446[0] = |(datain[311:308] ^ 11);
  assign w446[1] = |(datain[307:304] ^ 1);
  assign w446[2] = |(datain[303:300] ^ 0);
  assign w446[3] = |(datain[299:296] ^ 4);
  assign w446[4] = |(datain[295:292] ^ 13);
  assign w446[5] = |(datain[291:288] ^ 3);
  assign w446[6] = |(datain[287:284] ^ 14);
  assign w446[7] = |(datain[283:280] ^ 8);
  assign w446[8] = |(datain[279:276] ^ 8);
  assign w446[9] = |(datain[275:272] ^ 12);
  assign w446[10] = |(datain[271:268] ^ 13);
  assign w446[11] = |(datain[267:264] ^ 9);
  assign w446[12] = |(datain[263:260] ^ 0);
  assign w446[13] = |(datain[259:256] ^ 3);
  assign w446[14] = |(datain[255:252] ^ 12);
  assign w446[15] = |(datain[251:248] ^ 1);
  assign w446[16] = |(datain[247:244] ^ 11);
  assign w446[17] = |(datain[243:240] ^ 10);
  assign w446[18] = |(datain[239:236] ^ 0);
  assign w446[19] = |(datain[235:232] ^ 11);
  assign w446[20] = |(datain[231:228] ^ 0);
  assign w446[21] = |(datain[227:224] ^ 0);
  assign w446[22] = |(datain[223:220] ^ 14);
  assign w446[23] = |(datain[219:216] ^ 11);
  assign w446[24] = |(datain[215:212] ^ 7);
  assign w446[25] = |(datain[211:208] ^ 1);
  assign w446[26] = |(datain[207:204] ^ 11);
  assign w446[27] = |(datain[203:200] ^ 8);
  assign w446[28] = |(datain[199:196] ^ 13);
  assign w446[29] = |(datain[195:192] ^ 0);
  assign comp[446] = ~(|w446);
  wire [32-1:0] w447;
  assign w447[0] = |(datain[311:308] ^ 1);
  assign w447[1] = |(datain[307:304] ^ 15);
  assign w447[2] = |(datain[303:300] ^ 3);
  assign w447[3] = |(datain[299:296] ^ 2);
  assign w447[4] = |(datain[295:292] ^ 15);
  assign w447[5] = |(datain[291:288] ^ 6);
  assign w447[6] = |(datain[287:284] ^ 11);
  assign w447[7] = |(datain[283:280] ^ 9);
  assign w447[8] = |(datain[279:276] ^ 0);
  assign w447[9] = |(datain[275:272] ^ 2);
  assign w447[10] = |(datain[271:268] ^ 0);
  assign w447[11] = |(datain[267:264] ^ 0);
  assign w447[12] = |(datain[263:260] ^ 3);
  assign w447[13] = |(datain[259:256] ^ 3);
  assign w447[14] = |(datain[255:252] ^ 13);
  assign w447[15] = |(datain[251:248] ^ 11);
  assign w447[16] = |(datain[247:244] ^ 11);
  assign w447[17] = |(datain[243:240] ^ 8);
  assign w447[18] = |(datain[239:236] ^ 0);
  assign w447[19] = |(datain[235:232] ^ 2);
  assign w447[20] = |(datain[231:228] ^ 0);
  assign w447[21] = |(datain[227:224] ^ 2);
  assign w447[22] = |(datain[223:220] ^ 12);
  assign w447[23] = |(datain[219:216] ^ 13);
  assign w447[24] = |(datain[215:212] ^ 1);
  assign w447[25] = |(datain[211:208] ^ 3);
  assign w447[26] = |(datain[207:204] ^ 14);
  assign w447[27] = |(datain[203:200] ^ 9);
  assign w447[28] = |(datain[199:196] ^ 14);
  assign w447[29] = |(datain[195:192] ^ 14);
  assign w447[30] = |(datain[191:188] ^ 15);
  assign w447[31] = |(datain[187:184] ^ 14);
  assign comp[447] = ~(|w447);
  wire [42-1:0] w448;
  assign w448[0] = |(datain[311:308] ^ 11);
  assign w448[1] = |(datain[307:304] ^ 10);
  assign w448[2] = |(datain[303:300] ^ 2);
  assign w448[3] = |(datain[299:296] ^ 7);
  assign w448[4] = |(datain[295:292] ^ 0);
  assign w448[5] = |(datain[291:288] ^ 4);
  assign w448[6] = |(datain[287:284] ^ 5);
  assign w448[7] = |(datain[283:280] ^ 1);
  assign w448[8] = |(datain[279:276] ^ 5);
  assign w448[9] = |(datain[275:272] ^ 3);
  assign w448[10] = |(datain[271:268] ^ 5);
  assign w448[11] = |(datain[267:264] ^ 0);
  assign w448[12] = |(datain[263:260] ^ 5);
  assign w448[13] = |(datain[259:256] ^ 2);
  assign w448[14] = |(datain[255:252] ^ 12);
  assign w448[15] = |(datain[251:248] ^ 11);
  assign w448[16] = |(datain[247:244] ^ 8);
  assign w448[17] = |(datain[243:240] ^ 14);
  assign w448[18] = |(datain[239:236] ^ 12);
  assign w448[19] = |(datain[235:232] ^ 1);
  assign w448[20] = |(datain[231:228] ^ 11);
  assign w448[21] = |(datain[227:224] ^ 1);
  assign w448[22] = |(datain[223:220] ^ 0);
  assign w448[23] = |(datain[219:216] ^ 4);
  assign w448[24] = |(datain[215:212] ^ 11);
  assign w448[25] = |(datain[211:208] ^ 14);
  assign w448[26] = |(datain[207:204] ^ 11);
  assign w448[27] = |(datain[203:200] ^ 0);
  assign w448[28] = |(datain[199:196] ^ 0);
  assign w448[29] = |(datain[195:192] ^ 5);
  assign w448[30] = |(datain[191:188] ^ 8);
  assign w448[31] = |(datain[187:184] ^ 3);
  assign w448[32] = |(datain[183:180] ^ 12);
  assign w448[33] = |(datain[179:176] ^ 6);
  assign w448[34] = |(datain[175:172] ^ 0);
  assign w448[35] = |(datain[171:168] ^ 14);
  assign w448[36] = |(datain[167:164] ^ 10);
  assign w448[37] = |(datain[163:160] ^ 13);
  assign w448[38] = |(datain[159:156] ^ 3);
  assign w448[39] = |(datain[155:152] ^ 12);
  assign w448[40] = |(datain[151:148] ^ 8);
  assign w448[41] = |(datain[147:144] ^ 0);
  assign comp[448] = ~(|w448);
  wire [32-1:0] w449;
  assign w449[0] = |(datain[311:308] ^ 11);
  assign w449[1] = |(datain[307:304] ^ 4);
  assign w449[2] = |(datain[303:300] ^ 1);
  assign w449[3] = |(datain[299:296] ^ 3);
  assign w449[4] = |(datain[295:292] ^ 12);
  assign w449[5] = |(datain[291:288] ^ 13);
  assign w449[6] = |(datain[287:284] ^ 2);
  assign w449[7] = |(datain[283:280] ^ 15);
  assign w449[8] = |(datain[279:276] ^ 0);
  assign w449[9] = |(datain[275:272] ^ 6);
  assign w449[10] = |(datain[271:268] ^ 5);
  assign w449[11] = |(datain[267:264] ^ 3);
  assign w449[12] = |(datain[263:260] ^ 11);
  assign w449[13] = |(datain[259:256] ^ 4);
  assign w449[14] = |(datain[255:252] ^ 1);
  assign w449[15] = |(datain[251:248] ^ 3);
  assign w449[16] = |(datain[247:244] ^ 12);
  assign w449[17] = |(datain[243:240] ^ 13);
  assign w449[18] = |(datain[239:236] ^ 2);
  assign w449[19] = |(datain[235:232] ^ 15);
  assign w449[20] = |(datain[231:228] ^ 5);
  assign w449[21] = |(datain[227:224] ^ 8);
  assign w449[22] = |(datain[223:220] ^ 5);
  assign w449[23] = |(datain[219:216] ^ 10);
  assign w449[24] = |(datain[215:212] ^ 8);
  assign w449[25] = |(datain[211:208] ^ 7);
  assign w449[26] = |(datain[207:204] ^ 0);
  assign w449[27] = |(datain[203:200] ^ 4);
  assign w449[28] = |(datain[199:196] ^ 8);
  assign w449[29] = |(datain[195:192] ^ 7);
  assign w449[30] = |(datain[191:188] ^ 5);
  assign w449[31] = |(datain[187:184] ^ 4);
  assign comp[449] = ~(|w449);
  wire [28-1:0] w450;
  assign w450[0] = |(datain[311:308] ^ 12);
  assign w450[1] = |(datain[307:304] ^ 13);
  assign w450[2] = |(datain[303:300] ^ 2);
  assign w450[3] = |(datain[299:296] ^ 15);
  assign w450[4] = |(datain[295:292] ^ 5);
  assign w450[5] = |(datain[291:288] ^ 8);
  assign w450[6] = |(datain[287:284] ^ 5);
  assign w450[7] = |(datain[283:280] ^ 10);
  assign w450[8] = |(datain[279:276] ^ 8);
  assign w450[9] = |(datain[275:272] ^ 7);
  assign w450[10] = |(datain[271:268] ^ 0);
  assign w450[11] = |(datain[267:264] ^ 4);
  assign w450[12] = |(datain[263:260] ^ 8);
  assign w450[13] = |(datain[259:256] ^ 7);
  assign w450[14] = |(datain[255:252] ^ 5);
  assign w450[15] = |(datain[251:248] ^ 4);
  assign w450[16] = |(datain[247:244] ^ 0);
  assign w450[17] = |(datain[243:240] ^ 2);
  assign w450[18] = |(datain[239:236] ^ 5);
  assign w450[19] = |(datain[235:232] ^ 2);
  assign w450[20] = |(datain[231:228] ^ 5);
  assign w450[21] = |(datain[227:224] ^ 0);
  assign w450[22] = |(datain[223:220] ^ 5);
  assign w450[23] = |(datain[219:216] ^ 1);
  assign w450[24] = |(datain[215:212] ^ 5);
  assign w450[25] = |(datain[211:208] ^ 6);
  assign w450[26] = |(datain[207:204] ^ 10);
  assign w450[27] = |(datain[203:200] ^ 0);
  assign comp[450] = ~(|w450);
  wire [76-1:0] w451;
  assign w451[0] = |(datain[311:308] ^ 9);
  assign w451[1] = |(datain[307:304] ^ 7);
  assign w451[2] = |(datain[303:300] ^ 0);
  assign w451[3] = |(datain[299:296] ^ 3);
  assign w451[4] = |(datain[295:292] ^ 8);
  assign w451[5] = |(datain[291:288] ^ 9);
  assign w451[6] = |(datain[287:284] ^ 0);
  assign w451[7] = |(datain[283:280] ^ 13);
  assign w451[8] = |(datain[279:276] ^ 11);
  assign w451[9] = |(datain[275:272] ^ 9);
  assign w451[10] = |(datain[271:268] ^ 11);
  assign w451[11] = |(datain[267:264] ^ 6);
  assign w451[12] = |(datain[263:260] ^ 0);
  assign w451[13] = |(datain[259:256] ^ 3);
  assign w451[14] = |(datain[255:252] ^ 8);
  assign w451[15] = |(datain[251:248] ^ 11);
  assign w451[16] = |(datain[247:244] ^ 13);
  assign w451[17] = |(datain[243:240] ^ 6);
  assign w451[18] = |(datain[239:236] ^ 8);
  assign w451[19] = |(datain[235:232] ^ 1);
  assign w451[20] = |(datain[231:228] ^ 14);
  assign w451[21] = |(datain[227:224] ^ 10);
  assign w451[22] = |(datain[223:220] ^ 9);
  assign w451[23] = |(datain[219:216] ^ 12);
  assign w451[24] = |(datain[215:212] ^ 0);
  assign w451[25] = |(datain[211:208] ^ 3);
  assign w451[26] = |(datain[207:204] ^ 11);
  assign w451[27] = |(datain[203:200] ^ 4);
  assign w451[28] = |(datain[199:196] ^ 4);
  assign w451[29] = |(datain[195:192] ^ 0);
  assign w451[30] = |(datain[191:188] ^ 12);
  assign w451[31] = |(datain[187:184] ^ 13);
  assign w451[32] = |(datain[183:180] ^ 2);
  assign w451[33] = |(datain[179:176] ^ 1);
  assign w451[34] = |(datain[175:172] ^ 7);
  assign w451[35] = |(datain[171:168] ^ 2);
  assign w451[36] = |(datain[167:164] ^ 2);
  assign w451[37] = |(datain[163:160] ^ 1);
  assign w451[38] = |(datain[159:156] ^ 3);
  assign w451[39] = |(datain[155:152] ^ 3);
  assign w451[40] = |(datain[151:148] ^ 12);
  assign w451[41] = |(datain[147:144] ^ 9);
  assign w451[42] = |(datain[143:140] ^ 3);
  assign w451[43] = |(datain[139:136] ^ 3);
  assign w451[44] = |(datain[135:132] ^ 13);
  assign w451[45] = |(datain[131:128] ^ 2);
  assign w451[46] = |(datain[127:124] ^ 11);
  assign w451[47] = |(datain[123:120] ^ 8);
  assign w451[48] = |(datain[119:116] ^ 4);
  assign w451[49] = |(datain[115:112] ^ 2);
  assign w451[50] = |(datain[111:108] ^ 0);
  assign w451[51] = |(datain[107:104] ^ 0);
  assign w451[52] = |(datain[103:100] ^ 8);
  assign w451[53] = |(datain[99:96] ^ 6);
  assign w451[54] = |(datain[95:92] ^ 14);
  assign w451[55] = |(datain[91:88] ^ 0);
  assign w451[56] = |(datain[87:84] ^ 12);
  assign w451[57] = |(datain[83:80] ^ 13);
  assign w451[58] = |(datain[79:76] ^ 2);
  assign w451[59] = |(datain[75:72] ^ 1);
  assign w451[60] = |(datain[71:68] ^ 7);
  assign w451[61] = |(datain[67:64] ^ 2);
  assign w451[62] = |(datain[63:60] ^ 1);
  assign w451[63] = |(datain[59:56] ^ 4);
  assign w451[64] = |(datain[55:52] ^ 11);
  assign w451[65] = |(datain[51:48] ^ 9);
  assign w451[66] = |(datain[47:44] ^ 0);
  assign w451[67] = |(datain[43:40] ^ 3);
  assign w451[68] = |(datain[39:36] ^ 0);
  assign w451[69] = |(datain[35:32] ^ 0);
  assign w451[70] = |(datain[31:28] ^ 8);
  assign w451[71] = |(datain[27:24] ^ 1);
  assign w451[72] = |(datain[23:20] ^ 7);
  assign w451[73] = |(datain[19:16] ^ 12);
  assign w451[74] = |(datain[15:12] ^ 15);
  assign w451[75] = |(datain[11:8] ^ 14);
  assign comp[451] = ~(|w451);
  wire [46-1:0] w452;
  assign w452[0] = |(datain[311:308] ^ 8);
  assign w452[1] = |(datain[307:304] ^ 9);
  assign w452[2] = |(datain[303:300] ^ 4);
  assign w452[3] = |(datain[299:296] ^ 5);
  assign w452[4] = |(datain[295:292] ^ 1);
  assign w452[5] = |(datain[291:288] ^ 5);
  assign w452[6] = |(datain[287:284] ^ 11);
  assign w452[7] = |(datain[283:280] ^ 4);
  assign w452[8] = |(datain[279:276] ^ 4);
  assign w452[9] = |(datain[275:272] ^ 0);
  assign w452[10] = |(datain[271:268] ^ 11);
  assign w452[11] = |(datain[267:264] ^ 9);
  assign w452[12] = |(datain[263:260] ^ 13);
  assign w452[13] = |(datain[259:256] ^ 3);
  assign w452[14] = |(datain[255:252] ^ 0);
  assign w452[15] = |(datain[251:248] ^ 4);
  assign w452[16] = |(datain[247:244] ^ 11);
  assign w452[17] = |(datain[243:240] ^ 10);
  assign w452[18] = |(datain[239:236] ^ 0);
  assign w452[19] = |(datain[235:232] ^ 0);
  assign w452[20] = |(datain[231:228] ^ 0);
  assign w452[21] = |(datain[227:224] ^ 0);
  assign w452[22] = |(datain[223:220] ^ 12);
  assign w452[23] = |(datain[219:216] ^ 13);
  assign w452[24] = |(datain[215:212] ^ 2);
  assign w452[25] = |(datain[211:208] ^ 1);
  assign w452[26] = |(datain[207:204] ^ 11);
  assign w452[27] = |(datain[203:200] ^ 4);
  assign w452[28] = |(datain[199:196] ^ 3);
  assign w452[29] = |(datain[195:192] ^ 14);
  assign w452[30] = |(datain[191:188] ^ 12);
  assign w452[31] = |(datain[187:184] ^ 13);
  assign w452[32] = |(datain[183:180] ^ 2);
  assign w452[33] = |(datain[179:176] ^ 1);
  assign w452[34] = |(datain[175:172] ^ 5);
  assign w452[35] = |(datain[171:168] ^ 8);
  assign w452[36] = |(datain[167:164] ^ 2);
  assign w452[37] = |(datain[163:160] ^ 6);
  assign w452[38] = |(datain[159:156] ^ 8);
  assign w452[39] = |(datain[155:152] ^ 8);
  assign w452[40] = |(datain[151:148] ^ 4);
  assign w452[41] = |(datain[147:144] ^ 5);
  assign w452[42] = |(datain[143:140] ^ 0);
  assign w452[43] = |(datain[139:136] ^ 4);
  assign w452[44] = |(datain[135:132] ^ 14);
  assign w452[45] = |(datain[131:128] ^ 11);
  assign comp[452] = ~(|w452);
  wire [76-1:0] w453;
  assign w453[0] = |(datain[311:308] ^ 11);
  assign w453[1] = |(datain[307:304] ^ 14);
  assign w453[2] = |(datain[303:300] ^ 2);
  assign w453[3] = |(datain[299:296] ^ 9);
  assign w453[4] = |(datain[295:292] ^ 0);
  assign w453[5] = |(datain[291:288] ^ 1);
  assign w453[6] = |(datain[287:284] ^ 4);
  assign w453[7] = |(datain[283:280] ^ 1);
  assign w453[8] = |(datain[279:276] ^ 7);
  assign w453[9] = |(datain[275:272] ^ 4);
  assign w453[10] = |(datain[271:268] ^ 4);
  assign w453[11] = |(datain[267:264] ^ 1);
  assign w453[12] = |(datain[263:260] ^ 11);
  assign w453[13] = |(datain[259:256] ^ 8);
  assign w453[14] = |(datain[255:252] ^ 0);
  assign w453[15] = |(datain[251:248] ^ 2);
  assign w453[16] = |(datain[247:244] ^ 4);
  assign w453[17] = |(datain[243:240] ^ 2);
  assign w453[18] = |(datain[239:236] ^ 3);
  assign w453[19] = |(datain[235:232] ^ 3);
  assign w453[20] = |(datain[231:228] ^ 12);
  assign w453[21] = |(datain[227:224] ^ 9);
  assign w453[22] = |(datain[223:220] ^ 9);
  assign w453[23] = |(datain[219:216] ^ 9);
  assign w453[24] = |(datain[215:212] ^ 12);
  assign w453[25] = |(datain[211:208] ^ 13);
  assign w453[26] = |(datain[207:204] ^ 2);
  assign w453[27] = |(datain[203:200] ^ 1);
  assign w453[28] = |(datain[199:196] ^ 2);
  assign w453[29] = |(datain[195:192] ^ 13);
  assign w453[30] = |(datain[191:188] ^ 0);
  assign w453[31] = |(datain[187:184] ^ 3);
  assign w453[32] = |(datain[183:180] ^ 0);
  assign w453[33] = |(datain[179:176] ^ 0);
  assign w453[34] = |(datain[175:172] ^ 3);
  assign w453[35] = |(datain[171:168] ^ 14);
  assign w453[36] = |(datain[167:164] ^ 8);
  assign w453[37] = |(datain[163:160] ^ 9);
  assign w453[38] = |(datain[159:156] ^ 8);
  assign w453[39] = |(datain[155:152] ^ 6);
  assign w453[40] = |(datain[151:148] ^ 2);
  assign w453[41] = |(datain[147:144] ^ 11);
  assign w453[42] = |(datain[143:140] ^ 0);
  assign w453[43] = |(datain[139:136] ^ 1);
  assign w453[44] = |(datain[135:132] ^ 11);
  assign w453[45] = |(datain[131:128] ^ 4);
  assign w453[46] = |(datain[127:124] ^ 4);
  assign w453[47] = |(datain[123:120] ^ 0);
  assign w453[48] = |(datain[119:116] ^ 11);
  assign w453[49] = |(datain[115:112] ^ 9);
  assign w453[50] = |(datain[111:108] ^ 8);
  assign w453[51] = |(datain[107:104] ^ 5);
  assign w453[52] = |(datain[103:100] ^ 0);
  assign w453[53] = |(datain[99:96] ^ 3);
  assign w453[54] = |(datain[95:92] ^ 8);
  assign w453[55] = |(datain[91:88] ^ 13);
  assign w453[56] = |(datain[87:84] ^ 9);
  assign w453[57] = |(datain[83:80] ^ 6);
  assign w453[58] = |(datain[79:76] ^ 0);
  assign w453[59] = |(datain[75:72] ^ 0);
  assign w453[60] = |(datain[71:68] ^ 0);
  assign w453[61] = |(datain[67:64] ^ 1);
  assign w453[62] = |(datain[63:60] ^ 12);
  assign w453[63] = |(datain[59:56] ^ 13);
  assign w453[64] = |(datain[55:52] ^ 2);
  assign w453[65] = |(datain[51:48] ^ 1);
  assign w453[66] = |(datain[47:44] ^ 11);
  assign w453[67] = |(datain[43:40] ^ 8);
  assign w453[68] = |(datain[39:36] ^ 0);
  assign w453[69] = |(datain[35:32] ^ 0);
  assign w453[70] = |(datain[31:28] ^ 4);
  assign w453[71] = |(datain[27:24] ^ 2);
  assign w453[72] = |(datain[23:20] ^ 3);
  assign w453[73] = |(datain[19:16] ^ 3);
  assign w453[74] = |(datain[15:12] ^ 12);
  assign w453[75] = |(datain[11:8] ^ 9);
  assign comp[453] = ~(|w453);
  wire [46-1:0] w454;
  assign w454[0] = |(datain[311:308] ^ 0);
  assign w454[1] = |(datain[307:304] ^ 2);
  assign w454[2] = |(datain[303:300] ^ 4);
  assign w454[3] = |(datain[299:296] ^ 2);
  assign w454[4] = |(datain[295:292] ^ 9);
  assign w454[5] = |(datain[291:288] ^ 9);
  assign w454[6] = |(datain[287:284] ^ 3);
  assign w454[7] = |(datain[283:280] ^ 3);
  assign w454[8] = |(datain[279:276] ^ 12);
  assign w454[9] = |(datain[275:272] ^ 9);
  assign w454[10] = |(datain[271:268] ^ 12);
  assign w454[11] = |(datain[267:264] ^ 13);
  assign w454[12] = |(datain[263:260] ^ 2);
  assign w454[13] = |(datain[259:256] ^ 1);
  assign w454[14] = |(datain[255:252] ^ 11);
  assign w454[15] = |(datain[251:248] ^ 4);
  assign w454[16] = |(datain[247:244] ^ 4);
  assign w454[17] = |(datain[243:240] ^ 0);
  assign w454[18] = |(datain[239:236] ^ 8);
  assign w454[19] = |(datain[235:232] ^ 11);
  assign w454[20] = |(datain[231:228] ^ 13);
  assign w454[21] = |(datain[227:224] ^ 5);
  assign w454[22] = |(datain[223:220] ^ 11);
  assign w454[23] = |(datain[219:216] ^ 9);
  assign w454[24] = |(datain[215:212] ^ 11);
  assign w454[25] = |(datain[211:208] ^ 15);
  assign w454[26] = |(datain[207:204] ^ 0);
  assign w454[27] = |(datain[203:200] ^ 3);
  assign w454[28] = |(datain[199:196] ^ 12);
  assign w454[29] = |(datain[195:192] ^ 13);
  assign w454[30] = |(datain[191:188] ^ 2);
  assign w454[31] = |(datain[187:184] ^ 1);
  assign w454[32] = |(datain[183:180] ^ 11);
  assign w454[33] = |(datain[179:176] ^ 8);
  assign w454[34] = |(datain[175:172] ^ 0);
  assign w454[35] = |(datain[171:168] ^ 0);
  assign w454[36] = |(datain[167:164] ^ 4);
  assign w454[37] = |(datain[163:160] ^ 2);
  assign w454[38] = |(datain[159:156] ^ 9);
  assign w454[39] = |(datain[155:152] ^ 9);
  assign w454[40] = |(datain[151:148] ^ 3);
  assign w454[41] = |(datain[147:144] ^ 3);
  assign w454[42] = |(datain[143:140] ^ 12);
  assign w454[43] = |(datain[139:136] ^ 9);
  assign w454[44] = |(datain[135:132] ^ 12);
  assign w454[45] = |(datain[131:128] ^ 13);
  assign comp[454] = ~(|w454);
  wire [42-1:0] w455;
  assign w455[0] = |(datain[311:308] ^ 11);
  assign w455[1] = |(datain[307:304] ^ 10);
  assign w455[2] = |(datain[303:300] ^ 0);
  assign w455[3] = |(datain[299:296] ^ 0);
  assign w455[4] = |(datain[295:292] ^ 0);
  assign w455[5] = |(datain[291:288] ^ 1);
  assign w455[6] = |(datain[287:284] ^ 0);
  assign w455[7] = |(datain[283:280] ^ 14);
  assign w455[8] = |(datain[279:276] ^ 1);
  assign w455[9] = |(datain[275:272] ^ 15);
  assign w455[10] = |(datain[271:268] ^ 11);
  assign w455[11] = |(datain[267:264] ^ 4);
  assign w455[12] = |(datain[263:260] ^ 4);
  assign w455[13] = |(datain[259:256] ^ 0);
  assign w455[14] = |(datain[255:252] ^ 2);
  assign w455[15] = |(datain[251:248] ^ 14);
  assign w455[16] = |(datain[247:244] ^ 8);
  assign w455[17] = |(datain[243:240] ^ 11);
  assign w455[18] = |(datain[239:236] ^ 1);
  assign w455[19] = |(datain[235:232] ^ 14);
  assign w455[20] = |(datain[231:228] ^ 7);
  assign w455[21] = |(datain[227:224] ^ 0);
  assign w455[22] = |(datain[223:220] ^ 0);
  assign w455[23] = |(datain[219:216] ^ 3);
  assign w455[24] = |(datain[215:212] ^ 12);
  assign w455[25] = |(datain[211:208] ^ 13);
  assign w455[26] = |(datain[207:204] ^ 2);
  assign w455[27] = |(datain[203:200] ^ 1);
  assign w455[28] = |(datain[199:196] ^ 11);
  assign w455[29] = |(datain[195:192] ^ 8);
  assign w455[30] = |(datain[191:188] ^ 0);
  assign w455[31] = |(datain[187:184] ^ 2);
  assign w455[32] = |(datain[183:180] ^ 4);
  assign w455[33] = |(datain[179:176] ^ 2);
  assign w455[34] = |(datain[175:172] ^ 3);
  assign w455[35] = |(datain[171:168] ^ 3);
  assign w455[36] = |(datain[167:164] ^ 12);
  assign w455[37] = |(datain[163:160] ^ 9);
  assign w455[38] = |(datain[159:156] ^ 3);
  assign w455[39] = |(datain[155:152] ^ 3);
  assign w455[40] = |(datain[151:148] ^ 13);
  assign w455[41] = |(datain[147:144] ^ 2);
  assign comp[455] = ~(|w455);
  wire [76-1:0] w456;
  assign w456[0] = |(datain[311:308] ^ 5);
  assign w456[1] = |(datain[307:304] ^ 0);
  assign w456[2] = |(datain[303:300] ^ 5);
  assign w456[3] = |(datain[299:296] ^ 3);
  assign w456[4] = |(datain[295:292] ^ 8);
  assign w456[5] = |(datain[291:288] ^ 9);
  assign w456[6] = |(datain[287:284] ^ 2);
  assign w456[7] = |(datain[283:280] ^ 6);
  assign w456[8] = |(datain[279:276] ^ 5);
  assign w456[9] = |(datain[275:272] ^ 14);
  assign w456[10] = |(datain[271:268] ^ 0);
  assign w456[11] = |(datain[267:264] ^ 8);
  assign w456[12] = |(datain[263:260] ^ 8);
  assign w456[13] = |(datain[259:256] ^ 12);
  assign w456[14] = |(datain[255:252] ^ 1);
  assign w456[15] = |(datain[251:248] ^ 6);
  assign w456[16] = |(datain[247:244] ^ 6);
  assign w456[17] = |(datain[243:240] ^ 0);
  assign w456[18] = |(datain[239:236] ^ 0);
  assign w456[19] = |(datain[235:232] ^ 8);
  assign w456[20] = |(datain[231:228] ^ 0);
  assign w456[21] = |(datain[227:224] ^ 14);
  assign w456[22] = |(datain[223:220] ^ 1);
  assign w456[23] = |(datain[219:216] ^ 7);
  assign w456[24] = |(datain[215:212] ^ 11);
  assign w456[25] = |(datain[211:208] ^ 12);
  assign w456[26] = |(datain[207:204] ^ 0);
  assign w456[27] = |(datain[203:200] ^ 9);
  assign w456[28] = |(datain[199:196] ^ 0);
  assign w456[29] = |(datain[195:192] ^ 1);
  assign w456[30] = |(datain[191:188] ^ 2);
  assign w456[31] = |(datain[187:184] ^ 14);
  assign w456[32] = |(datain[183:180] ^ 10);
  assign w456[33] = |(datain[179:176] ^ 1);
  assign w456[34] = |(datain[175:172] ^ 0);
  assign w456[35] = |(datain[171:168] ^ 8);
  assign w456[36] = |(datain[167:164] ^ 0);
  assign w456[37] = |(datain[163:160] ^ 8);
  assign w456[38] = |(datain[159:156] ^ 5);
  assign w456[39] = |(datain[155:152] ^ 11);
  assign w456[40] = |(datain[151:148] ^ 3);
  assign w456[41] = |(datain[147:144] ^ 3);
  assign w456[42] = |(datain[143:140] ^ 13);
  assign w456[43] = |(datain[139:136] ^ 8);
  assign w456[44] = |(datain[135:132] ^ 5);
  assign w456[45] = |(datain[131:128] ^ 3);
  assign w456[46] = |(datain[127:124] ^ 5);
  assign w456[47] = |(datain[123:120] ^ 11);
  assign w456[48] = |(datain[119:116] ^ 8);
  assign w456[49] = |(datain[115:112] ^ 1);
  assign w456[50] = |(datain[111:108] ^ 15);
  assign w456[51] = |(datain[107:104] ^ 12);
  assign w456[52] = |(datain[103:100] ^ 0);
  assign w456[53] = |(datain[99:96] ^ 7);
  assign w456[54] = |(datain[95:92] ^ 0);
  assign w456[55] = |(datain[91:88] ^ 8);
  assign w456[56] = |(datain[87:84] ^ 7);
  assign w456[57] = |(datain[83:80] ^ 2);
  assign w456[58] = |(datain[79:76] ^ 15);
  assign w456[59] = |(datain[75:72] ^ 5);
  assign w456[60] = |(datain[71:68] ^ 8);
  assign w456[61] = |(datain[67:64] ^ 14);
  assign w456[62] = |(datain[63:60] ^ 1);
  assign w456[63] = |(datain[59:56] ^ 6);
  assign w456[64] = |(datain[55:52] ^ 6);
  assign w456[65] = |(datain[51:48] ^ 0);
  assign w456[66] = |(datain[47:44] ^ 0);
  assign w456[67] = |(datain[43:40] ^ 8);
  assign w456[68] = |(datain[39:36] ^ 8);
  assign w456[69] = |(datain[35:32] ^ 11);
  assign w456[70] = |(datain[31:28] ^ 2);
  assign w456[71] = |(datain[27:24] ^ 6);
  assign w456[72] = |(datain[23:20] ^ 5);
  assign w456[73] = |(datain[19:16] ^ 14);
  assign w456[74] = |(datain[15:12] ^ 0);
  assign w456[75] = |(datain[11:8] ^ 8);
  assign comp[456] = ~(|w456);
  wire [74-1:0] w457;
  assign w457[0] = |(datain[311:308] ^ 3);
  assign w457[1] = |(datain[307:304] ^ 3);
  assign w457[2] = |(datain[303:300] ^ 12);
  assign w457[3] = |(datain[299:296] ^ 9);
  assign w457[4] = |(datain[295:292] ^ 11);
  assign w457[5] = |(datain[291:288] ^ 8);
  assign w457[6] = |(datain[287:284] ^ 0);
  assign w457[7] = |(datain[283:280] ^ 1);
  assign w457[8] = |(datain[279:276] ^ 4);
  assign w457[9] = |(datain[275:272] ^ 3);
  assign w457[10] = |(datain[271:268] ^ 12);
  assign w457[11] = |(datain[267:264] ^ 13);
  assign w457[12] = |(datain[263:260] ^ 2);
  assign w457[13] = |(datain[259:256] ^ 1);
  assign w457[14] = |(datain[255:252] ^ 7);
  assign w457[15] = |(datain[251:248] ^ 2);
  assign w457[16] = |(datain[247:244] ^ 1);
  assign w457[17] = |(datain[243:240] ^ 9);
  assign w457[18] = |(datain[239:236] ^ 11);
  assign w457[19] = |(datain[235:232] ^ 8);
  assign w457[20] = |(datain[231:228] ^ 0);
  assign w457[21] = |(datain[227:224] ^ 1);
  assign w457[22] = |(datain[223:220] ^ 3);
  assign w457[23] = |(datain[219:216] ^ 13);
  assign w457[24] = |(datain[215:212] ^ 12);
  assign w457[25] = |(datain[211:208] ^ 13);
  assign w457[26] = |(datain[207:204] ^ 2);
  assign w457[27] = |(datain[203:200] ^ 1);
  assign w457[28] = |(datain[199:196] ^ 7);
  assign w457[29] = |(datain[195:192] ^ 2);
  assign w457[30] = |(datain[191:188] ^ 1);
  assign w457[31] = |(datain[187:184] ^ 2);
  assign w457[32] = |(datain[183:180] ^ 8);
  assign w457[33] = |(datain[179:176] ^ 11);
  assign w457[34] = |(datain[175:172] ^ 13);
  assign w457[35] = |(datain[171:168] ^ 8);
  assign w457[36] = |(datain[167:164] ^ 11);
  assign w457[37] = |(datain[163:160] ^ 10);
  assign w457[38] = |(datain[159:156] ^ 1);
  assign w457[39] = |(datain[155:152] ^ 6);
  assign w457[40] = |(datain[151:148] ^ 0);
  assign w457[41] = |(datain[147:144] ^ 2);
  assign w457[42] = |(datain[143:140] ^ 11);
  assign w457[43] = |(datain[139:136] ^ 4);
  assign w457[44] = |(datain[135:132] ^ 4);
  assign w457[45] = |(datain[131:128] ^ 0);
  assign w457[46] = |(datain[127:124] ^ 11);
  assign w457[47] = |(datain[123:120] ^ 9);
  assign w457[48] = |(datain[119:116] ^ 4);
  assign w457[49] = |(datain[115:112] ^ 9);
  assign w457[50] = |(datain[111:108] ^ 0);
  assign w457[51] = |(datain[107:104] ^ 0);
  assign w457[52] = |(datain[103:100] ^ 12);
  assign w457[53] = |(datain[99:96] ^ 13);
  assign w457[54] = |(datain[95:92] ^ 2);
  assign w457[55] = |(datain[91:88] ^ 1);
  assign w457[56] = |(datain[87:84] ^ 7);
  assign w457[57] = |(datain[83:80] ^ 2);
  assign w457[58] = |(datain[79:76] ^ 0);
  assign w457[59] = |(datain[75:72] ^ 4);
  assign w457[60] = |(datain[71:68] ^ 11);
  assign w457[61] = |(datain[67:64] ^ 4);
  assign w457[62] = |(datain[63:60] ^ 3);
  assign w457[63] = |(datain[59:56] ^ 14);
  assign w457[64] = |(datain[55:52] ^ 12);
  assign w457[65] = |(datain[51:48] ^ 13);
  assign w457[66] = |(datain[47:44] ^ 2);
  assign w457[67] = |(datain[43:40] ^ 1);
  assign w457[68] = |(datain[39:36] ^ 11);
  assign w457[69] = |(datain[35:32] ^ 10);
  assign w457[70] = |(datain[31:28] ^ 0);
  assign w457[71] = |(datain[27:24] ^ 0);
  assign w457[72] = |(datain[23:20] ^ 15);
  assign w457[73] = |(datain[19:16] ^ 15);
  assign comp[457] = ~(|w457);
  wire [76-1:0] w458;
  assign w458[0] = |(datain[311:308] ^ 10);
  assign w458[1] = |(datain[307:304] ^ 5);
  assign w458[2] = |(datain[303:300] ^ 0);
  assign w458[3] = |(datain[299:296] ^ 2);
  assign w458[4] = |(datain[295:292] ^ 11);
  assign w458[5] = |(datain[291:288] ^ 8);
  assign w458[6] = |(datain[287:284] ^ 0);
  assign w458[7] = |(datain[283:280] ^ 0);
  assign w458[8] = |(datain[279:276] ^ 10);
  assign w458[9] = |(datain[275:272] ^ 0);
  assign w458[10] = |(datain[271:268] ^ 8);
  assign w458[11] = |(datain[267:264] ^ 9);
  assign w458[12] = |(datain[263:260] ^ 8);
  assign w458[13] = |(datain[259:256] ^ 4);
  assign w458[14] = |(datain[255:252] ^ 9);
  assign w458[15] = |(datain[251:248] ^ 15);
  assign w458[16] = |(datain[247:244] ^ 0);
  assign w458[17] = |(datain[243:240] ^ 2);
  assign w458[18] = |(datain[239:236] ^ 11);
  assign w458[19] = |(datain[235:232] ^ 8);
  assign w458[20] = |(datain[231:228] ^ 0);
  assign w458[21] = |(datain[227:224] ^ 0);
  assign w458[22] = |(datain[223:220] ^ 4);
  assign w458[23] = |(datain[219:216] ^ 2);
  assign w458[24] = |(datain[215:212] ^ 3);
  assign w458[25] = |(datain[211:208] ^ 3);
  assign w458[26] = |(datain[207:204] ^ 12);
  assign w458[27] = |(datain[203:200] ^ 9);
  assign w458[28] = |(datain[199:196] ^ 3);
  assign w458[29] = |(datain[195:192] ^ 3);
  assign w458[30] = |(datain[191:188] ^ 13);
  assign w458[31] = |(datain[187:184] ^ 2);
  assign w458[32] = |(datain[183:180] ^ 12);
  assign w458[33] = |(datain[179:176] ^ 13);
  assign w458[34] = |(datain[175:172] ^ 3);
  assign w458[35] = |(datain[171:168] ^ 2);
  assign w458[36] = |(datain[167:164] ^ 11);
  assign w458[37] = |(datain[163:160] ^ 4);
  assign w458[38] = |(datain[159:156] ^ 4);
  assign w458[39] = |(datain[155:152] ^ 0);
  assign w458[40] = |(datain[151:148] ^ 11);
  assign w458[41] = |(datain[147:144] ^ 9);
  assign w458[42] = |(datain[143:140] ^ 1);
  assign w458[43] = |(datain[139:136] ^ 12);
  assign w458[44] = |(datain[135:132] ^ 0);
  assign w458[45] = |(datain[131:128] ^ 0);
  assign w458[46] = |(datain[127:124] ^ 11);
  assign w458[47] = |(datain[123:120] ^ 10);
  assign w458[48] = |(datain[119:116] ^ 8);
  assign w458[49] = |(datain[115:112] ^ 15);
  assign w458[50] = |(datain[111:108] ^ 0);
  assign w458[51] = |(datain[107:104] ^ 2);
  assign w458[52] = |(datain[103:100] ^ 0);
  assign w458[53] = |(datain[99:96] ^ 3);
  assign w458[54] = |(datain[95:92] ^ 13);
  assign w458[55] = |(datain[91:88] ^ 6);
  assign w458[56] = |(datain[87:84] ^ 12);
  assign w458[57] = |(datain[83:80] ^ 13);
  assign w458[58] = |(datain[79:76] ^ 3);
  assign w458[59] = |(datain[75:72] ^ 2);
  assign w458[60] = |(datain[71:68] ^ 7);
  assign w458[61] = |(datain[67:64] ^ 2);
  assign w458[62] = |(datain[63:60] ^ 2);
  assign w458[63] = |(datain[59:56] ^ 7);
  assign w458[64] = |(datain[55:52] ^ 5);
  assign w458[65] = |(datain[51:48] ^ 3);
  assign w458[66] = |(datain[47:44] ^ 11);
  assign w458[67] = |(datain[43:40] ^ 11);
  assign w458[68] = |(datain[39:36] ^ 6);
  assign w458[69] = |(datain[35:32] ^ 14);
  assign w458[70] = |(datain[31:28] ^ 0);
  assign w458[71] = |(datain[27:24] ^ 2);
  assign w458[72] = |(datain[23:20] ^ 0);
  assign w458[73] = |(datain[19:16] ^ 3);
  assign w458[74] = |(datain[15:12] ^ 13);
  assign w458[75] = |(datain[11:8] ^ 14);
  assign comp[458] = ~(|w458);
  wire [32-1:0] w459;
  assign w459[0] = |(datain[311:308] ^ 11);
  assign w459[1] = |(datain[307:304] ^ 8);
  assign w459[2] = |(datain[303:300] ^ 4);
  assign w459[3] = |(datain[299:296] ^ 0);
  assign w459[4] = |(datain[295:292] ^ 4);
  assign w459[5] = |(datain[291:288] ^ 11);
  assign w459[6] = |(datain[287:284] ^ 12);
  assign w459[7] = |(datain[283:280] ^ 13);
  assign w459[8] = |(datain[279:276] ^ 2);
  assign w459[9] = |(datain[275:272] ^ 1);
  assign w459[10] = |(datain[271:268] ^ 3);
  assign w459[11] = |(datain[267:264] ^ 13);
  assign w459[12] = |(datain[263:260] ^ 7);
  assign w459[13] = |(datain[259:256] ^ 8);
  assign w459[14] = |(datain[255:252] ^ 5);
  assign w459[15] = |(datain[251:248] ^ 6);
  assign w459[16] = |(datain[247:244] ^ 7);
  assign w459[17] = |(datain[243:240] ^ 5);
  assign w459[18] = |(datain[239:236] ^ 1);
  assign w459[19] = |(datain[235:232] ^ 2);
  assign w459[20] = |(datain[231:228] ^ 11);
  assign w459[21] = |(datain[227:224] ^ 8);
  assign w459[22] = |(datain[223:220] ^ 4);
  assign w459[23] = |(datain[219:216] ^ 1);
  assign w459[24] = |(datain[215:212] ^ 4);
  assign w459[25] = |(datain[211:208] ^ 11);
  assign w459[26] = |(datain[207:204] ^ 11);
  assign w459[27] = |(datain[203:200] ^ 15);
  assign w459[28] = |(datain[199:196] ^ 0);
  assign w459[29] = |(datain[195:192] ^ 0);
  assign w459[30] = |(datain[191:188] ^ 0);
  assign w459[31] = |(datain[187:184] ^ 1);
  assign comp[459] = ~(|w459);
  wire [38-1:0] w460;
  assign w460[0] = |(datain[311:308] ^ 1);
  assign w460[1] = |(datain[307:304] ^ 10);
  assign w460[2] = |(datain[303:300] ^ 0);
  assign w460[3] = |(datain[299:296] ^ 15);
  assign w460[4] = |(datain[295:292] ^ 5);
  assign w460[5] = |(datain[291:288] ^ 0);
  assign w460[6] = |(datain[287:284] ^ 12);
  assign w460[7] = |(datain[283:280] ^ 11);
  assign w460[8] = |(datain[279:276] ^ 2);
  assign w460[9] = |(datain[275:272] ^ 14);
  assign w460[10] = |(datain[271:268] ^ 8);
  assign w460[11] = |(datain[267:264] ^ 8);
  assign w460[12] = |(datain[263:260] ^ 1);
  assign w460[13] = |(datain[259:256] ^ 6);
  assign w460[14] = |(datain[255:252] ^ 4);
  assign w460[15] = |(datain[251:248] ^ 6);
  assign w460[16] = |(datain[247:244] ^ 0);
  assign w460[17] = |(datain[243:240] ^ 14);
  assign w460[18] = |(datain[239:236] ^ 3);
  assign w460[19] = |(datain[235:232] ^ 3);
  assign w460[20] = |(datain[231:228] ^ 12);
  assign w460[21] = |(datain[227:224] ^ 0);
  assign w460[22] = |(datain[223:220] ^ 8);
  assign w460[23] = |(datain[219:216] ^ 14);
  assign w460[24] = |(datain[215:212] ^ 13);
  assign w460[25] = |(datain[211:208] ^ 8);
  assign w460[26] = |(datain[207:204] ^ 12);
  assign w460[27] = |(datain[203:200] ^ 7);
  assign w460[28] = |(datain[199:196] ^ 0);
  assign w460[29] = |(datain[195:192] ^ 6);
  assign w460[30] = |(datain[191:188] ^ 8);
  assign w460[31] = |(datain[187:184] ^ 4);
  assign w460[32] = |(datain[183:180] ^ 0);
  assign w460[33] = |(datain[179:176] ^ 0);
  assign w460[34] = |(datain[175:172] ^ 15);
  assign w460[35] = |(datain[171:168] ^ 15);
  assign w460[36] = |(datain[167:164] ^ 15);
  assign w460[37] = |(datain[163:160] ^ 15);
  assign comp[460] = ~(|w460);
  wire [32-1:0] w461;
  assign w461[0] = |(datain[311:308] ^ 5);
  assign w461[1] = |(datain[307:304] ^ 9);
  assign w461[2] = |(datain[303:300] ^ 5);
  assign w461[3] = |(datain[299:296] ^ 11);
  assign w461[4] = |(datain[295:292] ^ 5);
  assign w461[5] = |(datain[291:288] ^ 8);
  assign w461[6] = |(datain[287:284] ^ 0);
  assign w461[7] = |(datain[283:280] ^ 7);
  assign w461[8] = |(datain[279:276] ^ 1);
  assign w461[9] = |(datain[275:272] ^ 15);
  assign w461[10] = |(datain[271:268] ^ 9);
  assign w461[11] = |(datain[267:264] ^ 12);
  assign w461[12] = |(datain[263:260] ^ 2);
  assign w461[13] = |(datain[259:256] ^ 14);
  assign w461[14] = |(datain[255:252] ^ 15);
  assign w461[15] = |(datain[251:248] ^ 15);
  assign w461[16] = |(datain[247:244] ^ 1);
  assign w461[17] = |(datain[243:240] ^ 14);
  assign w461[18] = |(datain[239:236] ^ 3);
  assign w461[19] = |(datain[235:232] ^ 11);
  assign w461[20] = |(datain[231:228] ^ 0);
  assign w461[21] = |(datain[227:224] ^ 0);
  assign w461[22] = |(datain[223:220] ^ 1);
  assign w461[23] = |(datain[219:216] ^ 14);
  assign w461[24] = |(datain[215:212] ^ 0);
  assign w461[25] = |(datain[211:208] ^ 7);
  assign w461[26] = |(datain[207:204] ^ 11);
  assign w461[27] = |(datain[203:200] ^ 4);
  assign w461[28] = |(datain[199:196] ^ 4);
  assign w461[29] = |(datain[195:192] ^ 9);
  assign w461[30] = |(datain[191:188] ^ 12);
  assign w461[31] = |(datain[187:184] ^ 13);
  assign comp[461] = ~(|w461);
  wire [30-1:0] w462;
  assign w462[0] = |(datain[311:308] ^ 8);
  assign w462[1] = |(datain[307:304] ^ 14);
  assign w462[2] = |(datain[303:300] ^ 13);
  assign w462[3] = |(datain[299:296] ^ 8);
  assign w462[4] = |(datain[295:292] ^ 10);
  assign w462[5] = |(datain[291:288] ^ 1);
  assign w462[6] = |(datain[287:284] ^ 1);
  assign w462[7] = |(datain[283:280] ^ 3);
  assign w462[8] = |(datain[279:276] ^ 0);
  assign w462[9] = |(datain[275:272] ^ 4);
  assign w462[10] = |(datain[271:268] ^ 11);
  assign w462[11] = |(datain[267:264] ^ 1);
  assign w462[12] = |(datain[263:260] ^ 0);
  assign w462[13] = |(datain[259:256] ^ 6);
  assign w462[14] = |(datain[255:252] ^ 13);
  assign w462[15] = |(datain[251:248] ^ 3);
  assign w462[16] = |(datain[247:244] ^ 14);
  assign w462[17] = |(datain[243:240] ^ 0);
  assign w462[18] = |(datain[239:236] ^ 8);
  assign w462[19] = |(datain[235:232] ^ 14);
  assign w462[20] = |(datain[231:228] ^ 13);
  assign w462[21] = |(datain[227:224] ^ 8);
  assign w462[22] = |(datain[223:220] ^ 3);
  assign w462[23] = |(datain[219:216] ^ 3);
  assign w462[24] = |(datain[215:212] ^ 15);
  assign w462[25] = |(datain[211:208] ^ 6);
  assign w462[26] = |(datain[207:204] ^ 8);
  assign w462[27] = |(datain[203:200] ^ 11);
  assign w462[28] = |(datain[199:196] ^ 4);
  assign w462[29] = |(datain[195:192] ^ 4);
  assign comp[462] = ~(|w462);
  wire [46-1:0] w463;
  assign w463[0] = |(datain[311:308] ^ 12);
  assign w463[1] = |(datain[307:304] ^ 0);
  assign w463[2] = |(datain[303:300] ^ 8);
  assign w463[3] = |(datain[299:296] ^ 14);
  assign w463[4] = |(datain[295:292] ^ 13);
  assign w463[5] = |(datain[291:288] ^ 8);
  assign w463[6] = |(datain[287:284] ^ 10);
  assign w463[7] = |(datain[283:280] ^ 0);
  assign w463[8] = |(datain[279:276] ^ 1);
  assign w463[9] = |(datain[275:272] ^ 7);
  assign w463[10] = |(datain[271:268] ^ 0);
  assign w463[11] = |(datain[267:264] ^ 4);
  assign w463[12] = |(datain[263:260] ^ 1);
  assign w463[13] = |(datain[259:256] ^ 15);
  assign w463[14] = |(datain[255:252] ^ 2);
  assign w463[15] = |(datain[251:248] ^ 4);
  assign w463[16] = |(datain[247:244] ^ 0);
  assign w463[17] = |(datain[243:240] ^ 12);
  assign w463[18] = |(datain[239:236] ^ 3);
  assign w463[19] = |(datain[235:232] ^ 12);
  assign w463[20] = |(datain[231:228] ^ 0);
  assign w463[21] = |(datain[227:224] ^ 12);
  assign w463[22] = |(datain[223:220] ^ 7);
  assign w463[23] = |(datain[219:216] ^ 5);
  assign w463[24] = |(datain[215:212] ^ 3);
  assign w463[25] = |(datain[211:208] ^ 4);
  assign w463[26] = |(datain[207:204] ^ 14);
  assign w463[27] = |(datain[203:200] ^ 4);
  assign w463[28] = |(datain[199:196] ^ 6);
  assign w463[29] = |(datain[195:192] ^ 0);
  assign w463[30] = |(datain[191:188] ^ 2);
  assign w463[31] = |(datain[187:184] ^ 4);
  assign w463[32] = |(datain[183:180] ^ 7);
  assign w463[33] = |(datain[179:176] ^ 15);
  assign w463[34] = |(datain[175:172] ^ 3);
  assign w463[35] = |(datain[171:168] ^ 12);
  assign w463[36] = |(datain[167:164] ^ 5);
  assign w463[37] = |(datain[163:160] ^ 3);
  assign w463[38] = |(datain[159:156] ^ 7);
  assign w463[39] = |(datain[155:152] ^ 5);
  assign w463[40] = |(datain[151:148] ^ 2);
  assign w463[41] = |(datain[147:144] ^ 12);
  assign w463[42] = |(datain[143:140] ^ 2);
  assign w463[43] = |(datain[139:136] ^ 14);
  assign w463[44] = |(datain[135:132] ^ 10);
  assign w463[45] = |(datain[131:128] ^ 1);
  assign comp[463] = ~(|w463);
  wire [76-1:0] w464;
  assign w464[0] = |(datain[311:308] ^ 12);
  assign w464[1] = |(datain[307:304] ^ 13);
  assign w464[2] = |(datain[303:300] ^ 1);
  assign w464[3] = |(datain[299:296] ^ 3);
  assign w464[4] = |(datain[295:292] ^ 7);
  assign w464[5] = |(datain[291:288] ^ 3);
  assign w464[6] = |(datain[287:284] ^ 0);
  assign w464[7] = |(datain[283:280] ^ 5);
  assign w464[8] = |(datain[279:276] ^ 8);
  assign w464[9] = |(datain[275:272] ^ 0);
  assign w464[10] = |(datain[271:268] ^ 14);
  assign w464[11] = |(datain[267:264] ^ 4);
  assign w464[12] = |(datain[263:260] ^ 12);
  assign w464[13] = |(datain[259:256] ^ 3);
  assign w464[14] = |(datain[255:252] ^ 7);
  assign w464[15] = |(datain[251:248] ^ 5);
  assign w464[16] = |(datain[247:244] ^ 0);
  assign w464[17] = |(datain[243:240] ^ 10);
  assign w464[18] = |(datain[239:236] ^ 15);
  assign w464[19] = |(datain[235:232] ^ 14);
  assign w464[20] = |(datain[231:228] ^ 12);
  assign w464[21] = |(datain[227:224] ^ 5);
  assign w464[22] = |(datain[223:220] ^ 3);
  assign w464[23] = |(datain[219:216] ^ 10);
  assign w464[24] = |(datain[215:212] ^ 2);
  assign w464[25] = |(datain[211:208] ^ 14);
  assign w464[26] = |(datain[207:204] ^ 4);
  assign w464[27] = |(datain[203:200] ^ 9);
  assign w464[28] = |(datain[199:196] ^ 0);
  assign w464[29] = |(datain[195:192] ^ 2);
  assign w464[30] = |(datain[191:188] ^ 7);
  assign w464[31] = |(datain[187:184] ^ 4);
  assign w464[32] = |(datain[183:180] ^ 0);
  assign w464[33] = |(datain[179:176] ^ 2);
  assign w464[34] = |(datain[175:172] ^ 14);
  assign w464[35] = |(datain[171:168] ^ 11);
  assign w464[36] = |(datain[167:164] ^ 14);
  assign w464[37] = |(datain[163:160] ^ 8);
  assign w464[38] = |(datain[159:156] ^ 12);
  assign w464[39] = |(datain[155:152] ^ 3);
  assign w464[40] = |(datain[151:148] ^ 11);
  assign w464[41] = |(datain[147:144] ^ 11);
  assign w464[42] = |(datain[143:140] ^ 0);
  assign w464[43] = |(datain[139:136] ^ 0);
  assign w464[44] = |(datain[135:132] ^ 0);
  assign w464[45] = |(datain[131:128] ^ 0);
  assign w464[46] = |(datain[127:124] ^ 12);
  assign w464[47] = |(datain[123:120] ^ 7);
  assign w464[48] = |(datain[119:116] ^ 0);
  assign w464[49] = |(datain[115:112] ^ 6);
  assign w464[50] = |(datain[111:108] ^ 4);
  assign w464[51] = |(datain[107:104] ^ 13);
  assign w464[52] = |(datain[103:100] ^ 0);
  assign w464[53] = |(datain[99:96] ^ 2);
  assign w464[54] = |(datain[95:92] ^ 0);
  assign w464[55] = |(datain[91:88] ^ 0);
  assign w464[56] = |(datain[87:84] ^ 0);
  assign w464[57] = |(datain[83:80] ^ 0);
  assign w464[58] = |(datain[79:76] ^ 10);
  assign w464[59] = |(datain[75:72] ^ 0);
  assign w464[60] = |(datain[71:68] ^ 4);
  assign w464[61] = |(datain[67:64] ^ 11);
  assign w464[62] = |(datain[63:60] ^ 0);
  assign w464[63] = |(datain[59:56] ^ 2);
  assign w464[64] = |(datain[55:52] ^ 11);
  assign w464[65] = |(datain[51:48] ^ 4);
  assign w464[66] = |(datain[47:44] ^ 0);
  assign w464[67] = |(datain[43:40] ^ 3);
  assign w464[68] = |(datain[39:36] ^ 12);
  assign w464[69] = |(datain[35:32] ^ 13);
  assign w464[70] = |(datain[31:28] ^ 1);
  assign w464[71] = |(datain[27:24] ^ 3);
  assign w464[72] = |(datain[23:20] ^ 15);
  assign w464[73] = |(datain[19:16] ^ 14);
  assign w464[74] = |(datain[15:12] ^ 12);
  assign w464[75] = |(datain[11:8] ^ 6);
  assign comp[464] = ~(|w464);
  wire [32-1:0] w465;
  assign w465[0] = |(datain[311:308] ^ 12);
  assign w465[1] = |(datain[307:304] ^ 0);
  assign w465[2] = |(datain[303:300] ^ 2);
  assign w465[3] = |(datain[299:296] ^ 14);
  assign w465[4] = |(datain[295:292] ^ 8);
  assign w465[5] = |(datain[291:288] ^ 11);
  assign w465[6] = |(datain[287:284] ^ 1);
  assign w465[7] = |(datain[283:280] ^ 6);
  assign w465[8] = |(datain[279:276] ^ 4);
  assign w465[9] = |(datain[275:272] ^ 6);
  assign w465[10] = |(datain[271:268] ^ 0);
  assign w465[11] = |(datain[267:264] ^ 14);
  assign w465[12] = |(datain[263:260] ^ 3);
  assign w465[13] = |(datain[259:256] ^ 3);
  assign w465[14] = |(datain[255:252] ^ 13);
  assign w465[15] = |(datain[251:248] ^ 11);
  assign w465[16] = |(datain[247:244] ^ 2);
  assign w465[17] = |(datain[243:240] ^ 14);
  assign w465[18] = |(datain[239:236] ^ 8);
  assign w465[19] = |(datain[235:232] ^ 11);
  assign w465[20] = |(datain[231:228] ^ 0);
  assign w465[21] = |(datain[227:224] ^ 14);
  assign w465[22] = |(datain[223:220] ^ 4);
  assign w465[23] = |(datain[219:216] ^ 4);
  assign w465[24] = |(datain[215:212] ^ 0);
  assign w465[25] = |(datain[211:208] ^ 14);
  assign w465[26] = |(datain[207:204] ^ 11);
  assign w465[27] = |(datain[203:200] ^ 8);
  assign w465[28] = |(datain[199:196] ^ 0);
  assign w465[29] = |(datain[195:192] ^ 8);
  assign w465[30] = |(datain[191:188] ^ 0);
  assign w465[31] = |(datain[187:184] ^ 2);
  assign comp[465] = ~(|w465);
  wire [32-1:0] w466;
  assign w466[0] = |(datain[311:308] ^ 11);
  assign w466[1] = |(datain[307:304] ^ 10);
  assign w466[2] = |(datain[303:300] ^ 2);
  assign w466[3] = |(datain[299:296] ^ 14);
  assign w466[4] = |(datain[295:292] ^ 0);
  assign w466[5] = |(datain[291:288] ^ 0);
  assign w466[6] = |(datain[287:284] ^ 11);
  assign w466[7] = |(datain[283:280] ^ 8);
  assign w466[8] = |(datain[279:276] ^ 0);
  assign w466[9] = |(datain[275:272] ^ 2);
  assign w466[10] = |(datain[271:268] ^ 3);
  assign w466[11] = |(datain[267:264] ^ 13);
  assign w466[12] = |(datain[263:260] ^ 12);
  assign w466[13] = |(datain[259:256] ^ 13);
  assign w466[14] = |(datain[255:252] ^ 2);
  assign w466[15] = |(datain[251:248] ^ 1);
  assign w466[16] = |(datain[247:244] ^ 11);
  assign w466[17] = |(datain[243:240] ^ 4);
  assign w466[18] = |(datain[239:236] ^ 4);
  assign w466[19] = |(datain[235:232] ^ 1);
  assign w466[20] = |(datain[231:228] ^ 12);
  assign w466[21] = |(datain[227:224] ^ 13);
  assign w466[22] = |(datain[223:220] ^ 2);
  assign w466[23] = |(datain[219:216] ^ 1);
  assign w466[24] = |(datain[215:212] ^ 8);
  assign w466[25] = |(datain[211:208] ^ 11);
  assign w466[26] = |(datain[207:204] ^ 4);
  assign w466[27] = |(datain[203:200] ^ 12);
  assign w466[28] = |(datain[199:196] ^ 1);
  assign w466[29] = |(datain[195:192] ^ 6);
  assign w466[30] = |(datain[191:188] ^ 0);
  assign w466[31] = |(datain[187:184] ^ 3);
  assign comp[466] = ~(|w466);
  wire [32-1:0] w467;
  assign w467[0] = |(datain[311:308] ^ 4);
  assign w467[1] = |(datain[307:304] ^ 12);
  assign w467[2] = |(datain[303:300] ^ 0);
  assign w467[3] = |(datain[299:296] ^ 0);
  assign w467[4] = |(datain[295:292] ^ 2);
  assign w467[5] = |(datain[291:288] ^ 14);
  assign w467[6] = |(datain[287:284] ^ 8);
  assign w467[7] = |(datain[283:280] ^ 9);
  assign w467[8] = |(datain[279:276] ^ 8);
  assign w467[9] = |(datain[275:272] ^ 4);
  assign w467[10] = |(datain[271:268] ^ 11);
  assign w467[11] = |(datain[267:264] ^ 13);
  assign w467[12] = |(datain[263:260] ^ 15);
  assign w467[13] = |(datain[259:256] ^ 13);
  assign w467[14] = |(datain[255:252] ^ 2);
  assign w467[15] = |(datain[251:248] ^ 14);
  assign w467[16] = |(datain[247:244] ^ 8);
  assign w467[17] = |(datain[243:240] ^ 12);
  assign w467[18] = |(datain[239:236] ^ 8);
  assign w467[19] = |(datain[235:232] ^ 4);
  assign w467[20] = |(datain[231:228] ^ 11);
  assign w467[21] = |(datain[227:224] ^ 15);
  assign w467[22] = |(datain[223:220] ^ 15);
  assign w467[23] = |(datain[219:216] ^ 13);
  assign w467[24] = |(datain[215:212] ^ 12);
  assign w467[25] = |(datain[211:208] ^ 4);
  assign w467[26] = |(datain[207:204] ^ 1);
  assign w467[27] = |(datain[203:200] ^ 14);
  assign w467[28] = |(datain[199:196] ^ 8);
  assign w467[29] = |(datain[195:192] ^ 4);
  assign w467[30] = |(datain[191:188] ^ 0);
  assign w467[31] = |(datain[187:184] ^ 0);
  assign comp[467] = ~(|w467);
  wire [30-1:0] w468;
  assign w468[0] = |(datain[311:308] ^ 8);
  assign w468[1] = |(datain[307:304] ^ 11);
  assign w468[2] = |(datain[303:300] ^ 8);
  assign w468[3] = |(datain[299:296] ^ 4);
  assign w468[4] = |(datain[295:292] ^ 8);
  assign w468[5] = |(datain[291:288] ^ 9);
  assign w468[6] = |(datain[287:284] ^ 15);
  assign w468[7] = |(datain[283:280] ^ 13);
  assign w468[8] = |(datain[279:276] ^ 2);
  assign w468[9] = |(datain[275:272] ^ 14);
  assign w468[10] = |(datain[271:268] ^ 10);
  assign w468[11] = |(datain[267:264] ^ 3);
  assign w468[12] = |(datain[263:260] ^ 0);
  assign w468[13] = |(datain[259:256] ^ 0);
  assign w468[14] = |(datain[255:252] ^ 0);
  assign w468[15] = |(datain[251:248] ^ 1);
  assign w468[16] = |(datain[247:244] ^ 2);
  assign w468[17] = |(datain[243:240] ^ 14);
  assign w468[18] = |(datain[239:236] ^ 8);
  assign w468[19] = |(datain[235:232] ^ 11);
  assign w468[20] = |(datain[231:228] ^ 8);
  assign w468[21] = |(datain[227:224] ^ 4);
  assign w468[22] = |(datain[223:220] ^ 8);
  assign w468[23] = |(datain[219:216] ^ 11);
  assign w468[24] = |(datain[215:212] ^ 15);
  assign w468[25] = |(datain[211:208] ^ 13);
  assign w468[26] = |(datain[207:204] ^ 2);
  assign w468[27] = |(datain[203:200] ^ 14);
  assign w468[28] = |(datain[199:196] ^ 10);
  assign w468[29] = |(datain[195:192] ^ 3);
  assign comp[468] = ~(|w468);
  wire [32-1:0] w469;
  assign w469[0] = |(datain[311:308] ^ 8);
  assign w469[1] = |(datain[307:304] ^ 6);
  assign w469[2] = |(datain[303:300] ^ 0);
  assign w469[3] = |(datain[299:296] ^ 0);
  assign w469[4] = |(datain[295:292] ^ 15);
  assign w469[5] = |(datain[291:288] ^ 11);
  assign w469[6] = |(datain[287:284] ^ 15);
  assign w469[7] = |(datain[283:280] ^ 14);
  assign w469[8] = |(datain[279:276] ^ 0);
  assign w469[9] = |(datain[275:272] ^ 14);
  assign w469[10] = |(datain[271:268] ^ 7);
  assign w469[11] = |(datain[267:264] ^ 11);
  assign w469[12] = |(datain[263:260] ^ 0);
  assign w469[13] = |(datain[259:256] ^ 4);
  assign w469[14] = |(datain[255:252] ^ 5);
  assign w469[15] = |(datain[251:248] ^ 14);
  assign w469[16] = |(datain[247:244] ^ 2);
  assign w469[17] = |(datain[243:240] ^ 14);
  assign w469[18] = |(datain[239:236] ^ 8);
  assign w469[19] = |(datain[235:232] ^ 1);
  assign w469[20] = |(datain[231:228] ^ 11);
  assign w469[21] = |(datain[227:224] ^ 12);
  assign w469[22] = |(datain[223:220] ^ 8);
  assign w469[23] = |(datain[219:216] ^ 9);
  assign w469[24] = |(datain[215:212] ^ 15);
  assign w469[25] = |(datain[211:208] ^ 13);
  assign w469[26] = |(datain[207:204] ^ 4);
  assign w469[27] = |(datain[203:200] ^ 13);
  assign w469[28] = |(datain[199:196] ^ 5);
  assign w469[29] = |(datain[195:192] ^ 10);
  assign w469[30] = |(datain[191:188] ^ 7);
  assign w469[31] = |(datain[187:184] ^ 5);
  assign comp[469] = ~(|w469);
  wire [50-1:0] w470;
  assign w470[0] = |(datain[311:308] ^ 12);
  assign w470[1] = |(datain[307:304] ^ 0);
  assign w470[2] = |(datain[303:300] ^ 8);
  assign w470[3] = |(datain[299:296] ^ 14);
  assign w470[4] = |(datain[295:292] ^ 12);
  assign w470[5] = |(datain[291:288] ^ 0);
  assign w470[6] = |(datain[287:284] ^ 12);
  assign w470[7] = |(datain[283:280] ^ 13);
  assign w470[8] = |(datain[279:276] ^ 1);
  assign w470[9] = |(datain[275:272] ^ 3);
  assign w470[10] = |(datain[271:268] ^ 0);
  assign w470[11] = |(datain[267:264] ^ 14);
  assign w470[12] = |(datain[263:260] ^ 1);
  assign w470[13] = |(datain[259:256] ^ 15);
  assign w470[14] = |(datain[255:252] ^ 8);
  assign w470[15] = |(datain[251:248] ^ 0);
  assign w470[16] = |(datain[247:244] ^ 3);
  assign w470[17] = |(datain[243:240] ^ 14);
  assign w470[18] = |(datain[239:236] ^ 0);
  assign w470[19] = |(datain[235:232] ^ 11);
  assign w470[20] = |(datain[231:228] ^ 0);
  assign w470[21] = |(datain[227:224] ^ 0);
  assign w470[22] = |(datain[223:220] ^ 0);
  assign w470[23] = |(datain[219:216] ^ 0);
  assign w470[24] = |(datain[215:212] ^ 7);
  assign w470[25] = |(datain[211:208] ^ 4);
  assign w470[26] = |(datain[207:204] ^ 2);
  assign w470[27] = |(datain[203:200] ^ 4);
  assign w470[28] = |(datain[199:196] ^ 11);
  assign w470[29] = |(datain[195:192] ^ 14);
  assign w470[30] = |(datain[191:188] ^ 10);
  assign w470[31] = |(datain[187:184] ^ 14);
  assign w470[32] = |(datain[183:180] ^ 0);
  assign w470[33] = |(datain[179:176] ^ 1);
  assign w470[34] = |(datain[175:172] ^ 8);
  assign w470[35] = |(datain[171:168] ^ 3);
  assign w470[36] = |(datain[167:164] ^ 12);
  assign w470[37] = |(datain[163:160] ^ 6);
  assign w470[38] = |(datain[159:156] ^ 1);
  assign w470[39] = |(datain[155:152] ^ 0);
  assign w470[40] = |(datain[151:148] ^ 8);
  assign w470[41] = |(datain[147:144] ^ 0);
  assign w470[42] = |(datain[143:140] ^ 3);
  assign w470[43] = |(datain[139:136] ^ 12);
  assign w470[44] = |(datain[135:132] ^ 8);
  assign w470[45] = |(datain[131:128] ^ 0);
  assign w470[46] = |(datain[127:124] ^ 7);
  assign w470[47] = |(datain[123:120] ^ 5);
  assign w470[48] = |(datain[119:116] ^ 15);
  assign w470[49] = |(datain[115:112] ^ 8);
  assign comp[470] = ~(|w470);
  wire [46-1:0] w471;
  assign w471[0] = |(datain[311:308] ^ 2);
  assign w471[1] = |(datain[307:304] ^ 6);
  assign w471[2] = |(datain[303:300] ^ 0);
  assign w471[3] = |(datain[299:296] ^ 3);
  assign w471[4] = |(datain[295:292] ^ 0);
  assign w471[5] = |(datain[291:288] ^ 0);
  assign w471[6] = |(datain[287:284] ^ 3);
  assign w471[7] = |(datain[283:280] ^ 13);
  assign w471[8] = |(datain[279:276] ^ 0);
  assign w471[9] = |(datain[275:272] ^ 2);
  assign w471[10] = |(datain[271:268] ^ 0);
  assign w471[11] = |(datain[267:264] ^ 0);
  assign w471[12] = |(datain[263:260] ^ 7);
  assign w471[13] = |(datain[259:256] ^ 3);
  assign w471[14] = |(datain[255:252] ^ 0);
  assign w471[15] = |(datain[251:248] ^ 3);
  assign w471[16] = |(datain[247:244] ^ 14);
  assign w471[17] = |(datain[243:240] ^ 8);
  assign w471[18] = |(datain[239:236] ^ 12);
  assign w471[19] = |(datain[235:232] ^ 12);
  assign w471[20] = |(datain[231:228] ^ 0);
  assign w471[21] = |(datain[227:224] ^ 0);
  assign w471[22] = |(datain[223:220] ^ 14);
  assign w471[23] = |(datain[219:216] ^ 8);
  assign w471[24] = |(datain[215:212] ^ 14);
  assign w471[25] = |(datain[211:208] ^ 8);
  assign w471[26] = |(datain[207:204] ^ 0);
  assign w471[27] = |(datain[203:200] ^ 0);
  assign w471[28] = |(datain[199:196] ^ 5);
  assign w471[29] = |(datain[195:192] ^ 8);
  assign w471[30] = |(datain[191:188] ^ 1);
  assign w471[31] = |(datain[187:184] ^ 15);
  assign w471[32] = |(datain[183:180] ^ 2);
  assign w471[33] = |(datain[179:176] ^ 14);
  assign w471[34] = |(datain[175:172] ^ 15);
  assign w471[35] = |(datain[171:168] ^ 15);
  assign w471[36] = |(datain[167:164] ^ 2);
  assign w471[37] = |(datain[163:160] ^ 14);
  assign w471[38] = |(datain[159:156] ^ 0);
  assign w471[39] = |(datain[155:152] ^ 7);
  assign w471[40] = |(datain[151:148] ^ 0);
  assign w471[41] = |(datain[147:144] ^ 0);
  assign w471[42] = |(datain[143:140] ^ 3);
  assign w471[43] = |(datain[139:136] ^ 3);
  assign w471[44] = |(datain[135:132] ^ 12);
  assign w471[45] = |(datain[131:128] ^ 0);
  assign comp[471] = ~(|w471);
  wire [76-1:0] w472;
  assign w472[0] = |(datain[311:308] ^ 11);
  assign w472[1] = |(datain[307:304] ^ 0);
  assign w472[2] = |(datain[303:300] ^ 6);
  assign w472[3] = |(datain[299:296] ^ 2);
  assign w472[4] = |(datain[295:292] ^ 14);
  assign w472[5] = |(datain[291:288] ^ 11);
  assign w472[6] = |(datain[287:284] ^ 15);
  assign w472[7] = |(datain[283:280] ^ 3);
  assign w472[8] = |(datain[279:276] ^ 10);
  assign w472[9] = |(datain[275:272] ^ 3);
  assign w472[10] = |(datain[271:268] ^ 1);
  assign w472[11] = |(datain[267:264] ^ 7);
  assign w472[12] = |(datain[263:260] ^ 0);
  assign w472[13] = |(datain[259:256] ^ 6);
  assign w472[14] = |(datain[255:252] ^ 11);
  assign w472[15] = |(datain[251:248] ^ 0);
  assign w472[16] = |(datain[247:244] ^ 0);
  assign w472[17] = |(datain[243:240] ^ 0);
  assign w472[18] = |(datain[239:236] ^ 10);
  assign w472[19] = |(datain[235:232] ^ 2);
  assign w472[20] = |(datain[231:228] ^ 6);
  assign w472[21] = |(datain[227:224] ^ 10);
  assign w472[22] = |(datain[223:220] ^ 0);
  assign w472[23] = |(datain[219:216] ^ 1);
  assign w472[24] = |(datain[215:212] ^ 11);
  assign w472[25] = |(datain[211:208] ^ 10);
  assign w472[26] = |(datain[207:204] ^ 6);
  assign w472[27] = |(datain[203:200] ^ 12);
  assign w472[28] = |(datain[199:196] ^ 0);
  assign w472[29] = |(datain[195:192] ^ 6);
  assign w472[30] = |(datain[191:188] ^ 8);
  assign w472[31] = |(datain[187:184] ^ 11);
  assign w472[32] = |(datain[183:180] ^ 1);
  assign w472[33] = |(datain[179:176] ^ 14);
  assign w472[34] = |(datain[175:172] ^ 6);
  assign w472[35] = |(datain[171:168] ^ 1);
  assign w472[36] = |(datain[167:164] ^ 0);
  assign w472[37] = |(datain[163:160] ^ 1);
  assign w472[38] = |(datain[159:156] ^ 10);
  assign w472[39] = |(datain[155:152] ^ 0);
  assign w472[40] = |(datain[151:148] ^ 6);
  assign w472[41] = |(datain[147:144] ^ 3);
  assign w472[42] = |(datain[143:140] ^ 0);
  assign w472[43] = |(datain[139:136] ^ 1);
  assign w472[44] = |(datain[135:132] ^ 11);
  assign w472[45] = |(datain[131:128] ^ 4);
  assign w472[46] = |(datain[127:124] ^ 4);
  assign w472[47] = |(datain[123:120] ^ 0);
  assign w472[48] = |(datain[119:116] ^ 2);
  assign w472[49] = |(datain[115:112] ^ 4);
  assign w472[50] = |(datain[111:108] ^ 0);
  assign w472[51] = |(datain[107:104] ^ 2);
  assign w472[52] = |(datain[103:100] ^ 3);
  assign w472[53] = |(datain[99:96] ^ 12);
  assign w472[54] = |(datain[95:92] ^ 0);
  assign w472[55] = |(datain[91:88] ^ 2);
  assign w472[56] = |(datain[87:84] ^ 7);
  assign w472[57] = |(datain[83:80] ^ 5);
  assign w472[58] = |(datain[79:76] ^ 1);
  assign w472[59] = |(datain[75:72] ^ 10);
  assign w472[60] = |(datain[71:68] ^ 3);
  assign w472[61] = |(datain[67:64] ^ 3);
  assign w472[62] = |(datain[63:60] ^ 12);
  assign w472[63] = |(datain[59:56] ^ 9);
  assign w472[64] = |(datain[55:52] ^ 5);
  assign w472[65] = |(datain[51:48] ^ 2);
  assign w472[66] = |(datain[47:44] ^ 5);
  assign w472[67] = |(datain[43:40] ^ 15);
  assign w472[68] = |(datain[39:36] ^ 8);
  assign w472[69] = |(datain[35:32] ^ 10);
  assign w472[70] = |(datain[31:28] ^ 0);
  assign w472[71] = |(datain[27:24] ^ 5);
  assign w472[72] = |(datain[23:20] ^ 3);
  assign w472[73] = |(datain[19:16] ^ 12);
  assign w472[74] = |(datain[15:12] ^ 0);
  assign w472[75] = |(datain[11:8] ^ 0);
  assign comp[472] = ~(|w472);
  wire [44-1:0] w473;
  assign w473[0] = |(datain[311:308] ^ 12);
  assign w473[1] = |(datain[307:304] ^ 6);
  assign w473[2] = |(datain[303:300] ^ 0);
  assign w473[3] = |(datain[299:296] ^ 6);
  assign w473[4] = |(datain[295:292] ^ 4);
  assign w473[5] = |(datain[291:288] ^ 8);
  assign w473[6] = |(datain[287:284] ^ 0);
  assign w473[7] = |(datain[283:280] ^ 1);
  assign w473[8] = |(datain[279:276] ^ 0);
  assign w473[9] = |(datain[275:272] ^ 0);
  assign w473[10] = |(datain[271:268] ^ 11);
  assign w473[11] = |(datain[267:264] ^ 4);
  assign w473[12] = |(datain[263:260] ^ 2);
  assign w473[13] = |(datain[259:256] ^ 10);
  assign w473[14] = |(datain[255:252] ^ 12);
  assign w473[15] = |(datain[251:248] ^ 13);
  assign w473[16] = |(datain[247:244] ^ 2);
  assign w473[17] = |(datain[243:240] ^ 1);
  assign w473[18] = |(datain[239:236] ^ 8);
  assign w473[19] = |(datain[235:232] ^ 1);
  assign w473[20] = |(datain[231:228] ^ 15);
  assign w473[21] = |(datain[227:224] ^ 9);
  assign w473[22] = |(datain[223:220] ^ 12);
  assign w473[23] = |(datain[219:216] ^ 4);
  assign w473[24] = |(datain[215:212] ^ 0);
  assign w473[25] = |(datain[211:208] ^ 7);
  assign w473[26] = |(datain[207:204] ^ 7);
  assign w473[27] = |(datain[203:200] ^ 2);
  assign w473[28] = |(datain[199:196] ^ 0);
  assign w473[29] = |(datain[195:192] ^ 12);
  assign w473[30] = |(datain[191:188] ^ 8);
  assign w473[31] = |(datain[187:184] ^ 1);
  assign w473[32] = |(datain[183:180] ^ 15);
  assign w473[33] = |(datain[179:176] ^ 10);
  assign w473[34] = |(datain[175:172] ^ 1);
  assign w473[35] = |(datain[171:168] ^ 1);
  assign w473[36] = |(datain[167:164] ^ 0);
  assign w473[37] = |(datain[163:160] ^ 8);
  assign w473[38] = |(datain[159:156] ^ 14);
  assign w473[39] = |(datain[155:152] ^ 11);
  assign w473[40] = |(datain[151:148] ^ 0);
  assign w473[41] = |(datain[147:144] ^ 6);
  assign w473[42] = |(datain[143:140] ^ 9);
  assign w473[43] = |(datain[139:136] ^ 0);
  assign comp[473] = ~(|w473);
  wire [28-1:0] w474;
  assign w474[0] = |(datain[311:308] ^ 12);
  assign w474[1] = |(datain[307:304] ^ 13);
  assign w474[2] = |(datain[303:300] ^ 2);
  assign w474[3] = |(datain[299:296] ^ 1);
  assign w474[4] = |(datain[295:292] ^ 11);
  assign w474[5] = |(datain[291:288] ^ 8);
  assign w474[6] = |(datain[287:284] ^ 0);
  assign w474[7] = |(datain[283:280] ^ 9);
  assign w474[8] = |(datain[279:276] ^ 3);
  assign w474[9] = |(datain[275:272] ^ 5);
  assign w474[10] = |(datain[271:268] ^ 12);
  assign w474[11] = |(datain[267:264] ^ 13);
  assign w474[12] = |(datain[263:260] ^ 2);
  assign w474[13] = |(datain[259:256] ^ 1);
  assign w474[14] = |(datain[255:252] ^ 8);
  assign w474[15] = |(datain[251:248] ^ 9);
  assign w474[16] = |(datain[247:244] ^ 1);
  assign w474[17] = |(datain[243:240] ^ 14);
  assign w474[18] = |(datain[239:236] ^ 4);
  assign w474[19] = |(datain[235:232] ^ 4);
  assign w474[20] = |(datain[231:228] ^ 0);
  assign w474[21] = |(datain[227:224] ^ 1);
  assign w474[22] = |(datain[223:220] ^ 8);
  assign w474[23] = |(datain[219:216] ^ 12);
  assign w474[24] = |(datain[215:212] ^ 0);
  assign w474[25] = |(datain[211:208] ^ 6);
  assign w474[26] = |(datain[207:204] ^ 4);
  assign w474[27] = |(datain[203:200] ^ 6);
  assign comp[474] = ~(|w474);
  wire [40-1:0] w475;
  assign w475[0] = |(datain[311:308] ^ 5);
  assign w475[1] = |(datain[307:304] ^ 13);
  assign w475[2] = |(datain[303:300] ^ 8);
  assign w475[3] = |(datain[299:296] ^ 1);
  assign w475[4] = |(datain[295:292] ^ 14);
  assign w475[5] = |(datain[291:288] ^ 13);
  assign w475[6] = |(datain[287:284] ^ 0);
  assign w475[7] = |(datain[283:280] ^ 9);
  assign w475[8] = |(datain[279:276] ^ 0);
  assign w475[9] = |(datain[275:272] ^ 1);
  assign w475[10] = |(datain[271:268] ^ 8);
  assign w475[11] = |(datain[267:264] ^ 13);
  assign w475[12] = |(datain[263:260] ^ 11);
  assign w475[13] = |(datain[259:256] ^ 6);
  assign w475[14] = |(datain[255:252] ^ 2);
  assign w475[15] = |(datain[251:248] ^ 3);
  assign w475[16] = |(datain[247:244] ^ 0);
  assign w475[17] = |(datain[243:240] ^ 1);
  assign w475[18] = |(datain[239:236] ^ 8);
  assign w475[19] = |(datain[235:232] ^ 11);
  assign w475[20] = |(datain[231:228] ^ 15);
  assign w475[21] = |(datain[227:224] ^ 14);
  assign w475[22] = |(datain[223:220] ^ 11);
  assign w475[23] = |(datain[219:216] ^ 9);
  assign w475[24] = |(datain[215:212] ^ 1);
  assign w475[25] = |(datain[211:208] ^ 4);
  assign w475[26] = |(datain[207:204] ^ 0);
  assign w475[27] = |(datain[203:200] ^ 2);
  assign w475[28] = |(datain[199:196] ^ 8);
  assign w475[29] = |(datain[195:192] ^ 10);
  assign w475[30] = |(datain[191:188] ^ 2);
  assign w475[31] = |(datain[187:184] ^ 6);
  assign w475[32] = |(datain[183:180] ^ 0);
  assign w475[33] = |(datain[179:176] ^ 5);
  assign w475[34] = |(datain[175:172] ^ 0);
  assign w475[35] = |(datain[171:168] ^ 1);
  assign w475[36] = |(datain[167:164] ^ 15);
  assign w475[37] = |(datain[163:160] ^ 14);
  assign w475[38] = |(datain[159:156] ^ 12);
  assign w475[39] = |(datain[155:152] ^ 12);
  assign comp[475] = ~(|w475);
  wire [76-1:0] w476;
  assign w476[0] = |(datain[311:308] ^ 9);
  assign w476[1] = |(datain[307:304] ^ 12);
  assign w476[2] = |(datain[303:300] ^ 5);
  assign w476[3] = |(datain[299:296] ^ 8);
  assign w476[4] = |(datain[295:292] ^ 15);
  assign w476[5] = |(datain[291:288] ^ 11);
  assign w476[6] = |(datain[287:284] ^ 10);
  assign w476[7] = |(datain[283:280] ^ 9);
  assign w476[8] = |(datain[279:276] ^ 0);
  assign w476[9] = |(datain[275:272] ^ 0);
  assign w476[10] = |(datain[271:268] ^ 2);
  assign w476[11] = |(datain[267:264] ^ 0);
  assign w476[12] = |(datain[263:260] ^ 0);
  assign w476[13] = |(datain[259:256] ^ 15);
  assign w476[14] = |(datain[255:252] ^ 8);
  assign w476[15] = |(datain[251:248] ^ 4);
  assign w476[16] = |(datain[247:244] ^ 9);
  assign w476[17] = |(datain[243:240] ^ 0);
  assign w476[18] = |(datain[239:236] ^ 0);
  assign w476[19] = |(datain[235:232] ^ 0);
  assign w476[20] = |(datain[231:228] ^ 6);
  assign w476[21] = |(datain[227:224] ^ 6);
  assign w476[22] = |(datain[223:220] ^ 11);
  assign w476[23] = |(datain[219:216] ^ 14);
  assign w476[24] = |(datain[215:212] ^ 4);
  assign w476[25] = |(datain[211:208] ^ 9);
  assign w476[26] = |(datain[207:204] ^ 5);
  assign w476[27] = |(datain[203:200] ^ 4);
  assign w476[28] = |(datain[199:196] ^ 4);
  assign w476[29] = |(datain[195:192] ^ 14);
  assign w476[30] = |(datain[191:188] ^ 4);
  assign w476[31] = |(datain[187:184] ^ 1);
  assign w476[32] = |(datain[183:180] ^ 11);
  assign w476[33] = |(datain[179:176] ^ 4);
  assign w476[34] = |(datain[175:172] ^ 3);
  assign w476[35] = |(datain[171:168] ^ 0);
  assign w476[36] = |(datain[167:164] ^ 12);
  assign w476[37] = |(datain[163:160] ^ 13);
  assign w476[38] = |(datain[159:156] ^ 2);
  assign w476[39] = |(datain[155:152] ^ 1);
  assign w476[40] = |(datain[151:148] ^ 6);
  assign w476[41] = |(datain[147:144] ^ 6);
  assign w476[42] = |(datain[143:140] ^ 8);
  assign w476[43] = |(datain[139:136] ^ 1);
  assign w476[44] = |(datain[135:132] ^ 15);
  assign w476[45] = |(datain[131:128] ^ 14);
  assign w476[46] = |(datain[127:124] ^ 2);
  assign w476[47] = |(datain[123:120] ^ 1);
  assign w476[48] = |(datain[119:116] ^ 4);
  assign w476[49] = |(datain[115:112] ^ 1);
  assign w476[50] = |(datain[111:108] ^ 5);
  assign w476[51] = |(datain[107:104] ^ 4);
  assign w476[52] = |(datain[103:100] ^ 4);
  assign w476[53] = |(datain[99:96] ^ 5);
  assign w476[54] = |(datain[95:92] ^ 7);
  assign w476[55] = |(datain[91:88] ^ 4);
  assign w476[56] = |(datain[87:84] ^ 7);
  assign w476[57] = |(datain[83:80] ^ 13);
  assign w476[58] = |(datain[79:76] ^ 9);
  assign w476[59] = |(datain[75:72] ^ 0);
  assign w476[60] = |(datain[71:68] ^ 9);
  assign w476[61] = |(datain[67:64] ^ 0);
  assign w476[62] = |(datain[63:60] ^ 3);
  assign w476[63] = |(datain[59:56] ^ 12);
  assign w476[64] = |(datain[55:52] ^ 0);
  assign w476[65] = |(datain[51:48] ^ 5);
  assign w476[66] = |(datain[47:44] ^ 7);
  assign w476[67] = |(datain[43:40] ^ 2);
  assign w476[68] = |(datain[39:36] ^ 7);
  assign w476[69] = |(datain[35:32] ^ 7);
  assign w476[70] = |(datain[31:28] ^ 9);
  assign w476[71] = |(datain[27:24] ^ 0);
  assign w476[72] = |(datain[23:20] ^ 9);
  assign w476[73] = |(datain[19:16] ^ 0);
  assign w476[74] = |(datain[15:12] ^ 11);
  assign w476[75] = |(datain[11:8] ^ 8);
  assign comp[476] = ~(|w476);
  wire [76-1:0] w477;
  assign w477[0] = |(datain[311:308] ^ 8);
  assign w477[1] = |(datain[307:304] ^ 14);
  assign w477[2] = |(datain[303:300] ^ 13);
  assign w477[3] = |(datain[299:296] ^ 15);
  assign w477[4] = |(datain[295:292] ^ 12);
  assign w477[5] = |(datain[291:288] ^ 4);
  assign w477[6] = |(datain[287:284] ^ 1);
  assign w477[7] = |(datain[283:280] ^ 6);
  assign w477[8] = |(datain[279:276] ^ 4);
  assign w477[9] = |(datain[275:272] ^ 12);
  assign w477[10] = |(datain[271:268] ^ 0);
  assign w477[11] = |(datain[267:264] ^ 0);
  assign w477[12] = |(datain[263:260] ^ 8);
  assign w477[13] = |(datain[259:256] ^ 9);
  assign w477[14] = |(datain[255:252] ^ 1);
  assign w477[15] = |(datain[251:248] ^ 6);
  assign w477[16] = |(datain[247:244] ^ 4);
  assign w477[17] = |(datain[243:240] ^ 12);
  assign w477[18] = |(datain[239:236] ^ 0);
  assign w477[19] = |(datain[235:232] ^ 3);
  assign w477[20] = |(datain[231:228] ^ 8);
  assign w477[21] = |(datain[227:224] ^ 12);
  assign w477[22] = |(datain[223:220] ^ 0);
  assign w477[23] = |(datain[219:216] ^ 6);
  assign w477[24] = |(datain[215:212] ^ 4);
  assign w477[25] = |(datain[211:208] ^ 14);
  assign w477[26] = |(datain[207:204] ^ 0);
  assign w477[27] = |(datain[203:200] ^ 3);
  assign w477[28] = |(datain[199:196] ^ 15);
  assign w477[29] = |(datain[195:192] ^ 10);
  assign w477[30] = |(datain[191:188] ^ 8);
  assign w477[31] = |(datain[187:184] ^ 14);
  assign w477[32] = |(datain[183:180] ^ 13);
  assign w477[33] = |(datain[179:176] ^ 7);
  assign w477[34] = |(datain[175:172] ^ 11);
  assign w477[35] = |(datain[171:168] ^ 14);
  assign w477[36] = |(datain[167:164] ^ 0);
  assign w477[37] = |(datain[163:160] ^ 0);
  assign w477[38] = |(datain[159:156] ^ 7);
  assign w477[39] = |(datain[155:152] ^ 12);
  assign w477[40] = |(datain[151:148] ^ 8);
  assign w477[41] = |(datain[147:144] ^ 11);
  assign w477[42] = |(datain[143:140] ^ 14);
  assign w477[43] = |(datain[139:136] ^ 6);
  assign w477[44] = |(datain[135:132] ^ 15);
  assign w477[45] = |(datain[131:128] ^ 11);
  assign w477[46] = |(datain[127:124] ^ 1);
  assign w477[47] = |(datain[123:120] ^ 14);
  assign w477[48] = |(datain[119:116] ^ 5);
  assign w477[49] = |(datain[115:112] ^ 6);
  assign w477[50] = |(datain[111:108] ^ 5);
  assign w477[51] = |(datain[107:104] ^ 6);
  assign w477[52] = |(datain[103:100] ^ 10);
  assign w477[53] = |(datain[99:96] ^ 1);
  assign w477[54] = |(datain[95:92] ^ 1);
  assign w477[55] = |(datain[91:88] ^ 3);
  assign w477[56] = |(datain[87:84] ^ 0);
  assign w477[57] = |(datain[83:80] ^ 4);
  assign w477[58] = |(datain[79:76] ^ 4);
  assign w477[59] = |(datain[75:72] ^ 8);
  assign w477[60] = |(datain[71:68] ^ 10);
  assign w477[61] = |(datain[67:64] ^ 3);
  assign w477[62] = |(datain[63:60] ^ 1);
  assign w477[63] = |(datain[59:56] ^ 3);
  assign w477[64] = |(datain[55:52] ^ 0);
  assign w477[65] = |(datain[51:48] ^ 4);
  assign w477[66] = |(datain[47:44] ^ 11);
  assign w477[67] = |(datain[43:40] ^ 1);
  assign w477[68] = |(datain[39:36] ^ 0);
  assign w477[69] = |(datain[35:32] ^ 6);
  assign w477[70] = |(datain[31:28] ^ 13);
  assign w477[71] = |(datain[27:24] ^ 3);
  assign w477[72] = |(datain[23:20] ^ 14);
  assign w477[73] = |(datain[19:16] ^ 0);
  assign w477[74] = |(datain[15:12] ^ 8);
  assign w477[75] = |(datain[11:8] ^ 14);
  assign comp[477] = ~(|w477);
  wire [28-1:0] w478;
  assign w478[0] = |(datain[311:308] ^ 7);
  assign w478[1] = |(datain[307:304] ^ 4);
  assign w478[2] = |(datain[303:300] ^ 0);
  assign w478[3] = |(datain[299:296] ^ 15);
  assign w478[4] = |(datain[295:292] ^ 8);
  assign w478[5] = |(datain[291:288] ^ 0);
  assign w478[6] = |(datain[287:284] ^ 3);
  assign w478[7] = |(datain[283:280] ^ 14);
  assign w478[8] = |(datain[279:276] ^ 13);
  assign w478[9] = |(datain[275:272] ^ 14);
  assign w478[10] = |(datain[271:268] ^ 0);
  assign w478[11] = |(datain[267:264] ^ 3);
  assign w478[12] = |(datain[263:260] ^ 0);
  assign w478[13] = |(datain[259:256] ^ 2);
  assign w478[14] = |(datain[255:252] ^ 7);
  assign w478[15] = |(datain[251:248] ^ 4);
  assign w478[16] = |(datain[247:244] ^ 0);
  assign w478[17] = |(datain[243:240] ^ 12);
  assign w478[18] = |(datain[239:236] ^ 8);
  assign w478[19] = |(datain[235:232] ^ 0);
  assign w478[20] = |(datain[231:228] ^ 3);
  assign w478[21] = |(datain[227:224] ^ 14);
  assign w478[22] = |(datain[223:220] ^ 13);
  assign w478[23] = |(datain[219:216] ^ 14);
  assign w478[24] = |(datain[215:212] ^ 0);
  assign w478[25] = |(datain[211:208] ^ 3);
  assign w478[26] = |(datain[207:204] ^ 0);
  assign w478[27] = |(datain[203:200] ^ 3);
  assign comp[478] = ~(|w478);
  wire [70-1:0] w479;
  assign w479[0] = |(datain[311:308] ^ 0);
  assign w479[1] = |(datain[307:304] ^ 5);
  assign w479[2] = |(datain[303:300] ^ 0);
  assign w479[3] = |(datain[299:296] ^ 2);
  assign w479[4] = |(datain[295:292] ^ 0);
  assign w479[5] = |(datain[291:288] ^ 0);
  assign w479[6] = |(datain[287:284] ^ 5);
  assign w479[7] = |(datain[283:280] ^ 0);
  assign w479[8] = |(datain[279:276] ^ 12);
  assign w479[9] = |(datain[275:272] ^ 10);
  assign w479[10] = |(datain[271:268] ^ 0);
  assign w479[11] = |(datain[267:264] ^ 2);
  assign w479[12] = |(datain[263:260] ^ 0);
  assign w479[13] = |(datain[259:256] ^ 0);
  assign w479[14] = |(datain[255:252] ^ 5);
  assign w479[15] = |(datain[251:248] ^ 11);
  assign w479[16] = |(datain[247:244] ^ 8);
  assign w479[17] = |(datain[243:240] ^ 13);
  assign w479[18] = |(datain[239:236] ^ 5);
  assign w479[19] = |(datain[235:232] ^ 7);
  assign w479[20] = |(datain[231:228] ^ 0);
  assign w479[21] = |(datain[227:224] ^ 5);
  assign w479[22] = |(datain[223:220] ^ 2);
  assign w479[23] = |(datain[219:216] ^ 14);
  assign w479[24] = |(datain[215:212] ^ 8);
  assign w479[25] = |(datain[211:208] ^ 9);
  assign w479[26] = |(datain[207:204] ^ 1);
  assign w479[27] = |(datain[203:200] ^ 7);
  assign w479[28] = |(datain[199:196] ^ 2);
  assign w479[29] = |(datain[195:192] ^ 14);
  assign w479[30] = |(datain[191:188] ^ 8);
  assign w479[31] = |(datain[187:184] ^ 12);
  assign w479[32] = |(datain[183:180] ^ 4);
  assign w479[33] = |(datain[179:176] ^ 15);
  assign w479[34] = |(datain[175:172] ^ 0);
  assign w479[35] = |(datain[171:168] ^ 2);
  assign w479[36] = |(datain[167:164] ^ 9);
  assign w479[37] = |(datain[163:160] ^ 12);
  assign w479[38] = |(datain[159:156] ^ 2);
  assign w479[39] = |(datain[155:152] ^ 14);
  assign w479[40] = |(datain[151:148] ^ 15);
  assign w479[41] = |(datain[147:144] ^ 15);
  assign w479[42] = |(datain[143:140] ^ 1);
  assign w479[43] = |(datain[139:136] ^ 15);
  assign w479[44] = |(datain[135:132] ^ 12);
  assign w479[45] = |(datain[131:128] ^ 3);
  assign w479[46] = |(datain[127:124] ^ 0);
  assign w479[47] = |(datain[123:120] ^ 0);
  assign w479[48] = |(datain[119:116] ^ 2);
  assign w479[49] = |(datain[115:112] ^ 14);
  assign w479[50] = |(datain[111:108] ^ 8);
  assign w479[51] = |(datain[107:104] ^ 9);
  assign w479[52] = |(datain[103:100] ^ 2);
  assign w479[53] = |(datain[99:96] ^ 7);
  assign w479[54] = |(datain[95:92] ^ 8);
  assign w479[55] = |(datain[91:88] ^ 3);
  assign w479[56] = |(datain[87:84] ^ 12);
  assign w479[57] = |(datain[83:80] ^ 3);
  assign w479[58] = |(datain[79:76] ^ 2);
  assign w479[59] = |(datain[75:72] ^ 12);
  assign w479[60] = |(datain[71:68] ^ 8);
  assign w479[61] = |(datain[67:64] ^ 11);
  assign w479[62] = |(datain[63:60] ^ 14);
  assign w479[63] = |(datain[59:56] ^ 3);
  assign w479[64] = |(datain[55:52] ^ 5);
  assign w479[65] = |(datain[51:48] ^ 8);
  assign w479[66] = |(datain[47:44] ^ 5);
  assign w479[67] = |(datain[43:40] ^ 8);
  assign w479[68] = |(datain[39:36] ^ 3);
  assign w479[69] = |(datain[35:32] ^ 5);
  assign comp[479] = ~(|w479);
  wire [46-1:0] w480;
  assign w480[0] = |(datain[311:308] ^ 11);
  assign w480[1] = |(datain[307:304] ^ 15);
  assign w480[2] = |(datain[303:300] ^ 0);
  assign w480[3] = |(datain[299:296] ^ 5);
  assign w480[4] = |(datain[295:292] ^ 0);
  assign w480[5] = |(datain[291:288] ^ 6);
  assign w480[6] = |(datain[287:284] ^ 15);
  assign w480[7] = |(datain[283:280] ^ 12);
  assign w480[8] = |(datain[279:276] ^ 11);
  assign w480[9] = |(datain[275:272] ^ 0);
  assign w480[10] = |(datain[271:268] ^ 13);
  assign w480[11] = |(datain[267:264] ^ 9);
  assign w480[12] = |(datain[263:260] ^ 11);
  assign w480[13] = |(datain[259:256] ^ 14);
  assign w480[14] = |(datain[255:252] ^ 1);
  assign w480[15] = |(datain[251:248] ^ 9);
  assign w480[16] = |(datain[247:244] ^ 0);
  assign w480[17] = |(datain[243:240] ^ 0);
  assign w480[18] = |(datain[239:236] ^ 9);
  assign w480[19] = |(datain[235:232] ^ 0);
  assign w480[20] = |(datain[231:228] ^ 2);
  assign w480[21] = |(datain[227:224] ^ 14);
  assign w480[22] = |(datain[223:220] ^ 3);
  assign w480[23] = |(datain[219:216] ^ 0);
  assign w480[24] = |(datain[215:212] ^ 0);
  assign w480[25] = |(datain[211:208] ^ 4);
  assign w480[26] = |(datain[207:204] ^ 9);
  assign w480[27] = |(datain[203:200] ^ 0);
  assign w480[28] = |(datain[199:196] ^ 9);
  assign w480[29] = |(datain[195:192] ^ 0);
  assign w480[30] = |(datain[191:188] ^ 4);
  assign w480[31] = |(datain[187:184] ^ 6);
  assign w480[32] = |(datain[183:180] ^ 4);
  assign w480[33] = |(datain[179:176] ^ 15);
  assign w480[34] = |(datain[175:172] ^ 9);
  assign w480[35] = |(datain[171:168] ^ 0);
  assign w480[36] = |(datain[167:164] ^ 7);
  assign w480[37] = |(datain[163:160] ^ 5);
  assign w480[38] = |(datain[159:156] ^ 15);
  assign w480[39] = |(datain[155:152] ^ 5);
  assign w480[40] = |(datain[151:148] ^ 15);
  assign w480[41] = |(datain[147:144] ^ 12);
  assign w480[42] = |(datain[143:140] ^ 14);
  assign w480[43] = |(datain[139:136] ^ 11);
  assign w480[44] = |(datain[135:132] ^ 0);
  assign w480[45] = |(datain[131:128] ^ 0);
  assign comp[480] = ~(|w480);
  wire [44-1:0] w481;
  assign w481[0] = |(datain[311:308] ^ 0);
  assign w481[1] = |(datain[307:304] ^ 1);
  assign w481[2] = |(datain[303:300] ^ 8);
  assign w481[3] = |(datain[299:296] ^ 10);
  assign w481[4] = |(datain[295:292] ^ 2);
  assign w481[5] = |(datain[291:288] ^ 6);
  assign w481[6] = |(datain[287:284] ^ 0);
  assign w481[7] = |(datain[283:280] ^ 5);
  assign w481[8] = |(datain[279:276] ^ 0);
  assign w481[9] = |(datain[275:272] ^ 1);
  assign w481[10] = |(datain[271:268] ^ 14);
  assign w481[11] = |(datain[267:264] ^ 11);
  assign w481[12] = |(datain[263:260] ^ 1);
  assign w481[13] = |(datain[259:256] ^ 1);
  assign w481[14] = |(datain[255:252] ^ 10);
  assign w481[15] = |(datain[251:248] ^ 12);
  assign w481[16] = |(datain[247:244] ^ 3);
  assign w481[17] = |(datain[243:240] ^ 2);
  assign w481[18] = |(datain[239:236] ^ 12);
  assign w481[19] = |(datain[235:232] ^ 4);
  assign w481[20] = |(datain[231:228] ^ 10);
  assign w481[21] = |(datain[227:224] ^ 10);
  assign w481[22] = |(datain[223:220] ^ 14);
  assign w481[23] = |(datain[219:216] ^ 2);
  assign w481[24] = |(datain[215:212] ^ 15);
  assign w481[25] = |(datain[211:208] ^ 10);
  assign w481[26] = |(datain[207:204] ^ 11);
  assign w481[27] = |(datain[203:200] ^ 4);
  assign w481[28] = |(datain[199:196] ^ 1);
  assign w481[29] = |(datain[195:192] ^ 9);
  assign w481[30] = |(datain[191:188] ^ 12);
  assign w481[31] = |(datain[187:184] ^ 13);
  assign w481[32] = |(datain[183:180] ^ 2);
  assign w481[33] = |(datain[179:176] ^ 1);
  assign w481[34] = |(datain[175:172] ^ 8);
  assign w481[35] = |(datain[171:168] ^ 10);
  assign w481[36] = |(datain[167:164] ^ 15);
  assign w481[37] = |(datain[163:160] ^ 0);
  assign w481[38] = |(datain[159:156] ^ 11);
  assign w481[39] = |(datain[155:152] ^ 4);
  assign w481[40] = |(datain[151:148] ^ 0);
  assign w481[41] = |(datain[147:144] ^ 14);
  assign w481[42] = |(datain[143:140] ^ 12);
  assign w481[43] = |(datain[139:136] ^ 13);
  assign comp[481] = ~(|w481);
  wire [42-1:0] w482;
  assign w482[0] = |(datain[311:308] ^ 8);
  assign w482[1] = |(datain[307:304] ^ 10);
  assign w482[2] = |(datain[303:300] ^ 2);
  assign w482[3] = |(datain[299:296] ^ 6);
  assign w482[4] = |(datain[295:292] ^ 0);
  assign w482[5] = |(datain[291:288] ^ 7);
  assign w482[6] = |(datain[287:284] ^ 0);
  assign w482[7] = |(datain[283:280] ^ 1);
  assign w482[8] = |(datain[279:276] ^ 14);
  assign w482[9] = |(datain[275:272] ^ 11);
  assign w482[10] = |(datain[271:268] ^ 1);
  assign w482[11] = |(datain[267:264] ^ 2);
  assign w482[12] = |(datain[263:260] ^ 9);
  assign w482[13] = |(datain[259:256] ^ 0);
  assign w482[14] = |(datain[255:252] ^ 10);
  assign w482[15] = |(datain[251:248] ^ 12);
  assign w482[16] = |(datain[247:244] ^ 3);
  assign w482[17] = |(datain[243:240] ^ 2);
  assign w482[18] = |(datain[239:236] ^ 12);
  assign w482[19] = |(datain[235:232] ^ 4);
  assign w482[20] = |(datain[231:228] ^ 10);
  assign w482[21] = |(datain[227:224] ^ 10);
  assign w482[22] = |(datain[223:220] ^ 14);
  assign w482[23] = |(datain[219:216] ^ 2);
  assign w482[24] = |(datain[215:212] ^ 15);
  assign w482[25] = |(datain[211:208] ^ 10);
  assign w482[26] = |(datain[207:204] ^ 11);
  assign w482[27] = |(datain[203:200] ^ 4);
  assign w482[28] = |(datain[199:196] ^ 1);
  assign w482[29] = |(datain[195:192] ^ 9);
  assign w482[30] = |(datain[191:188] ^ 12);
  assign w482[31] = |(datain[187:184] ^ 13);
  assign w482[32] = |(datain[183:180] ^ 2);
  assign w482[33] = |(datain[179:176] ^ 1);
  assign w482[34] = |(datain[175:172] ^ 8);
  assign w482[35] = |(datain[171:168] ^ 10);
  assign w482[36] = |(datain[167:164] ^ 15);
  assign w482[37] = |(datain[163:160] ^ 0);
  assign w482[38] = |(datain[159:156] ^ 11);
  assign w482[39] = |(datain[155:152] ^ 4);
  assign w482[40] = |(datain[151:148] ^ 0);
  assign w482[41] = |(datain[147:144] ^ 14);
  assign comp[482] = ~(|w482);
  wire [30-1:0] w483;
  assign w483[0] = |(datain[311:308] ^ 5);
  assign w483[1] = |(datain[307:304] ^ 0);
  assign w483[2] = |(datain[303:300] ^ 5);
  assign w483[3] = |(datain[299:296] ^ 2);
  assign w483[4] = |(datain[295:292] ^ 11);
  assign w483[5] = |(datain[291:288] ^ 4);
  assign w483[6] = |(datain[287:284] ^ 1);
  assign w483[7] = |(datain[283:280] ^ 9);
  assign w483[8] = |(datain[279:276] ^ 12);
  assign w483[9] = |(datain[275:272] ^ 13);
  assign w483[10] = |(datain[271:268] ^ 2);
  assign w483[11] = |(datain[267:264] ^ 1);
  assign w483[12] = |(datain[263:260] ^ 8);
  assign w483[13] = |(datain[259:256] ^ 10);
  assign w483[14] = |(datain[255:252] ^ 13);
  assign w483[15] = |(datain[251:248] ^ 0);
  assign w483[16] = |(datain[247:244] ^ 11);
  assign w483[17] = |(datain[243:240] ^ 4);
  assign w483[18] = |(datain[239:236] ^ 0);
  assign w483[19] = |(datain[235:232] ^ 14);
  assign w483[20] = |(datain[231:228] ^ 12);
  assign w483[21] = |(datain[227:224] ^ 13);
  assign w483[22] = |(datain[223:220] ^ 2);
  assign w483[23] = |(datain[219:216] ^ 1);
  assign w483[24] = |(datain[215:212] ^ 3);
  assign w483[25] = |(datain[211:208] ^ 12);
  assign w483[26] = |(datain[207:204] ^ 0);
  assign w483[27] = |(datain[203:200] ^ 4);
  assign w483[28] = |(datain[199:196] ^ 7);
  assign w483[29] = |(datain[195:192] ^ 2);
  assign comp[483] = ~(|w483);
  wire [36-1:0] w484;
  assign w484[0] = |(datain[311:308] ^ 0);
  assign w484[1] = |(datain[307:304] ^ 6);
  assign w484[2] = |(datain[303:300] ^ 0);
  assign w484[3] = |(datain[299:296] ^ 2);
  assign w484[4] = |(datain[295:292] ^ 7);
  assign w484[5] = |(datain[291:288] ^ 2);
  assign w484[6] = |(datain[287:284] ^ 2);
  assign w484[7] = |(datain[283:280] ^ 14);
  assign w484[8] = |(datain[279:276] ^ 14);
  assign w484[9] = |(datain[275:272] ^ 8);
  assign w484[10] = |(datain[271:268] ^ 9);
  assign w484[11] = |(datain[267:264] ^ 1);
  assign w484[12] = |(datain[263:260] ^ 0);
  assign w484[13] = |(datain[259:256] ^ 0);
  assign w484[14] = |(datain[255:252] ^ 8);
  assign w484[15] = |(datain[251:248] ^ 13);
  assign w484[16] = |(datain[247:244] ^ 1);
  assign w484[17] = |(datain[243:240] ^ 6);
  assign w484[18] = |(datain[239:236] ^ 7);
  assign w484[19] = |(datain[235:232] ^ 2);
  assign w484[20] = |(datain[231:228] ^ 0);
  assign w484[21] = |(datain[227:224] ^ 5);
  assign w484[22] = |(datain[223:220] ^ 14);
  assign w484[23] = |(datain[219:216] ^ 8);
  assign w484[24] = |(datain[215:212] ^ 9);
  assign w484[25] = |(datain[211:208] ^ 7);
  assign w484[26] = |(datain[207:204] ^ 0);
  assign w484[27] = |(datain[203:200] ^ 0);
  assign w484[28] = |(datain[199:196] ^ 14);
  assign w484[29] = |(datain[195:192] ^ 8);
  assign w484[30] = |(datain[191:188] ^ 2);
  assign w484[31] = |(datain[187:184] ^ 3);
  assign w484[32] = |(datain[183:180] ^ 0);
  assign w484[33] = |(datain[179:176] ^ 0);
  assign w484[34] = |(datain[175:172] ^ 14);
  assign w484[35] = |(datain[171:168] ^ 8);
  assign comp[484] = ~(|w484);
  wire [42-1:0] w485;
  assign w485[0] = |(datain[311:308] ^ 2);
  assign w485[1] = |(datain[307:304] ^ 11);
  assign w485[2] = |(datain[303:300] ^ 13);
  assign w485[3] = |(datain[299:296] ^ 0);
  assign w485[4] = |(datain[295:292] ^ 3);
  assign w485[5] = |(datain[291:288] ^ 3);
  assign w485[6] = |(datain[287:284] ^ 12);
  assign w485[7] = |(datain[283:280] ^ 9);
  assign w485[8] = |(datain[279:276] ^ 11);
  assign w485[9] = |(datain[275:272] ^ 8);
  assign w485[10] = |(datain[271:268] ^ 0);
  assign w485[11] = |(datain[267:264] ^ 0);
  assign w485[12] = |(datain[263:260] ^ 4);
  assign w485[13] = |(datain[259:256] ^ 2);
  assign w485[14] = |(datain[255:252] ^ 12);
  assign w485[15] = |(datain[251:248] ^ 13);
  assign w485[16] = |(datain[247:244] ^ 2);
  assign w485[17] = |(datain[243:240] ^ 1);
  assign w485[18] = |(datain[239:236] ^ 11);
  assign w485[19] = |(datain[235:232] ^ 10);
  assign w485[20] = |(datain[231:228] ^ 0);
  assign w485[21] = |(datain[227:224] ^ 0);
  assign w485[22] = |(datain[223:220] ^ 0);
  assign w485[23] = |(datain[219:216] ^ 1);
  assign w485[24] = |(datain[215:212] ^ 11);
  assign w485[25] = |(datain[211:208] ^ 9);
  assign w485[26] = |(datain[207:204] ^ 10);
  assign w485[27] = |(datain[203:200] ^ 10);
  assign w485[28] = |(datain[199:196] ^ 0);
  assign w485[29] = |(datain[195:192] ^ 5);
  assign w485[30] = |(datain[191:188] ^ 11);
  assign w485[31] = |(datain[187:184] ^ 4);
  assign w485[32] = |(datain[183:180] ^ 4);
  assign w485[33] = |(datain[179:176] ^ 0);
  assign w485[34] = |(datain[175:172] ^ 12);
  assign w485[35] = |(datain[171:168] ^ 13);
  assign w485[36] = |(datain[167:164] ^ 2);
  assign w485[37] = |(datain[163:160] ^ 1);
  assign w485[38] = |(datain[159:156] ^ 5);
  assign w485[39] = |(datain[155:152] ^ 10);
  assign w485[40] = |(datain[151:148] ^ 5);
  assign w485[41] = |(datain[147:144] ^ 9);
  assign comp[485] = ~(|w485);
  wire [72-1:0] w486;
  assign w486[0] = |(datain[311:308] ^ 0);
  assign w486[1] = |(datain[307:304] ^ 1);
  assign w486[2] = |(datain[303:300] ^ 11);
  assign w486[3] = |(datain[299:296] ^ 4);
  assign w486[4] = |(datain[295:292] ^ 3);
  assign w486[5] = |(datain[291:288] ^ 14);
  assign w486[6] = |(datain[287:284] ^ 12);
  assign w486[7] = |(datain[283:280] ^ 13);
  assign w486[8] = |(datain[279:276] ^ 2);
  assign w486[9] = |(datain[275:272] ^ 1);
  assign w486[10] = |(datain[271:268] ^ 7);
  assign w486[11] = |(datain[267:264] ^ 2);
  assign w486[12] = |(datain[263:260] ^ 10);
  assign w486[13] = |(datain[259:256] ^ 5);
  assign w486[14] = |(datain[255:252] ^ 11);
  assign w486[15] = |(datain[251:248] ^ 4);
  assign w486[16] = |(datain[247:244] ^ 3);
  assign w486[17] = |(datain[243:240] ^ 12);
  assign w486[18] = |(datain[239:236] ^ 11);
  assign w486[19] = |(datain[235:232] ^ 9);
  assign w486[20] = |(datain[231:228] ^ 0);
  assign w486[21] = |(datain[227:224] ^ 0);
  assign w486[22] = |(datain[223:220] ^ 0);
  assign w486[23] = |(datain[219:216] ^ 0);
  assign w486[24] = |(datain[215:212] ^ 11);
  assign w486[25] = |(datain[211:208] ^ 10);
  assign w486[26] = |(datain[207:204] ^ 0);
  assign w486[27] = |(datain[203:200] ^ 3);
  assign w486[28] = |(datain[199:196] ^ 0);
  assign w486[29] = |(datain[195:192] ^ 1);
  assign w486[30] = |(datain[191:188] ^ 12);
  assign w486[31] = |(datain[187:184] ^ 13);
  assign w486[32] = |(datain[183:180] ^ 2);
  assign w486[33] = |(datain[179:176] ^ 1);
  assign w486[34] = |(datain[175:172] ^ 7);
  assign w486[35] = |(datain[171:168] ^ 2);
  assign w486[36] = |(datain[167:164] ^ 9);
  assign w486[37] = |(datain[163:160] ^ 9);
  assign w486[38] = |(datain[159:156] ^ 10);
  assign w486[39] = |(datain[155:152] ^ 3);
  assign w486[40] = |(datain[151:148] ^ 2);
  assign w486[41] = |(datain[147:144] ^ 5);
  assign w486[42] = |(datain[143:140] ^ 0);
  assign w486[43] = |(datain[139:136] ^ 1);
  assign w486[44] = |(datain[135:132] ^ 0);
  assign w486[45] = |(datain[131:128] ^ 6);
  assign w486[46] = |(datain[127:124] ^ 8);
  assign w486[47] = |(datain[123:120] ^ 11);
  assign w486[48] = |(datain[119:116] ^ 1);
  assign w486[49] = |(datain[115:112] ^ 14);
  assign w486[50] = |(datain[111:108] ^ 2);
  assign w486[51] = |(datain[107:104] ^ 9);
  assign w486[52] = |(datain[103:100] ^ 0);
  assign w486[53] = |(datain[99:96] ^ 1);
  assign w486[54] = |(datain[95:92] ^ 5);
  assign w486[55] = |(datain[91:88] ^ 3);
  assign w486[56] = |(datain[87:84] ^ 0);
  assign w486[57] = |(datain[83:80] ^ 7);
  assign w486[58] = |(datain[79:76] ^ 11);
  assign w486[59] = |(datain[75:72] ^ 9);
  assign w486[60] = |(datain[71:68] ^ 1);
  assign w486[61] = |(datain[67:64] ^ 14);
  assign w486[62] = |(datain[63:60] ^ 0);
  assign w486[63] = |(datain[59:56] ^ 0);
  assign w486[64] = |(datain[55:52] ^ 8);
  assign w486[65] = |(datain[51:48] ^ 11);
  assign w486[66] = |(datain[47:44] ^ 3);
  assign w486[67] = |(datain[43:40] ^ 6);
  assign w486[68] = |(datain[39:36] ^ 9);
  assign w486[69] = |(datain[35:32] ^ 1);
  assign w486[70] = |(datain[31:28] ^ 0);
  assign w486[71] = |(datain[27:24] ^ 1);
  assign comp[486] = ~(|w486);
  wire [46-1:0] w487;
  assign w487[0] = |(datain[311:308] ^ 11);
  assign w487[1] = |(datain[307:304] ^ 8);
  assign w487[2] = |(datain[303:300] ^ 0);
  assign w487[3] = |(datain[299:296] ^ 1);
  assign w487[4] = |(datain[295:292] ^ 9);
  assign w487[5] = |(datain[291:288] ^ 0);
  assign w487[6] = |(datain[287:284] ^ 8);
  assign w487[7] = |(datain[283:280] ^ 13);
  assign w487[8] = |(datain[279:276] ^ 9);
  assign w487[9] = |(datain[275:272] ^ 4);
  assign w487[10] = |(datain[271:268] ^ 0);
  assign w487[11] = |(datain[267:264] ^ 6);
  assign w487[12] = |(datain[263:260] ^ 0);
  assign w487[13] = |(datain[259:256] ^ 1);
  assign w487[14] = |(datain[255:252] ^ 11);
  assign w487[15] = |(datain[251:248] ^ 4);
  assign w487[16] = |(datain[247:244] ^ 4);
  assign w487[17] = |(datain[243:240] ^ 0);
  assign w487[18] = |(datain[239:236] ^ 12);
  assign w487[19] = |(datain[235:232] ^ 13);
  assign w487[20] = |(datain[231:228] ^ 2);
  assign w487[21] = |(datain[227:224] ^ 1);
  assign w487[22] = |(datain[223:220] ^ 7);
  assign w487[23] = |(datain[219:216] ^ 2);
  assign w487[24] = |(datain[215:212] ^ 2);
  assign w487[25] = |(datain[211:208] ^ 2);
  assign w487[26] = |(datain[207:204] ^ 5);
  assign w487[27] = |(datain[203:200] ^ 8);
  assign w487[28] = |(datain[199:196] ^ 0);
  assign w487[29] = |(datain[195:192] ^ 5);
  assign w487[30] = |(datain[191:188] ^ 5);
  assign w487[31] = |(datain[187:184] ^ 2);
  assign w487[32] = |(datain[183:180] ^ 0);
  assign w487[33] = |(datain[179:176] ^ 0);
  assign w487[34] = |(datain[175:172] ^ 12);
  assign w487[35] = |(datain[171:168] ^ 6);
  assign w487[36] = |(datain[167:164] ^ 0);
  assign w487[37] = |(datain[163:160] ^ 5);
  assign w487[38] = |(datain[159:156] ^ 14);
  assign w487[39] = |(datain[155:152] ^ 9);
  assign w487[40] = |(datain[151:148] ^ 8);
  assign w487[41] = |(datain[147:144] ^ 9);
  assign w487[42] = |(datain[143:140] ^ 4);
  assign w487[43] = |(datain[139:136] ^ 5);
  assign w487[44] = |(datain[135:132] ^ 0);
  assign w487[45] = |(datain[131:128] ^ 1);
  assign comp[487] = ~(|w487);
  wire [32-1:0] w488;
  assign w488[0] = |(datain[311:308] ^ 14);
  assign w488[1] = |(datain[307:304] ^ 8);
  assign w488[2] = |(datain[303:300] ^ 0);
  assign w488[3] = |(datain[299:296] ^ 0);
  assign w488[4] = |(datain[295:292] ^ 0);
  assign w488[5] = |(datain[291:288] ^ 0);
  assign w488[6] = |(datain[287:284] ^ 5);
  assign w488[7] = |(datain[283:280] ^ 14);
  assign w488[8] = |(datain[279:276] ^ 8);
  assign w488[9] = |(datain[275:272] ^ 1);
  assign w488[10] = |(datain[271:268] ^ 14);
  assign w488[11] = |(datain[267:264] ^ 14);
  assign w488[12] = |(datain[263:260] ^ 6);
  assign w488[13] = |(datain[259:256] ^ 5);
  assign w488[14] = |(datain[255:252] ^ 0);
  assign w488[15] = |(datain[251:248] ^ 1);
  assign w488[16] = |(datain[247:244] ^ 8);
  assign w488[17] = |(datain[243:240] ^ 8);
  assign w488[18] = |(datain[239:236] ^ 8);
  assign w488[19] = |(datain[235:232] ^ 4);
  assign w488[20] = |(datain[231:228] ^ 5);
  assign w488[21] = |(datain[227:224] ^ 4);
  assign w488[22] = |(datain[223:220] ^ 0);
  assign w488[23] = |(datain[219:216] ^ 1);
  assign w488[24] = |(datain[215:212] ^ 8);
  assign w488[25] = |(datain[211:208] ^ 11);
  assign w488[26] = |(datain[207:204] ^ 8);
  assign w488[27] = |(datain[203:200] ^ 4);
  assign w488[28] = |(datain[199:196] ^ 0);
  assign w488[29] = |(datain[195:192] ^ 6);
  assign w488[30] = |(datain[191:188] ^ 0);
  assign w488[31] = |(datain[187:184] ^ 1);
  assign comp[488] = ~(|w488);
  wire [20-1:0] w489;
  assign w489[0] = |(datain[311:308] ^ 5);
  assign w489[1] = |(datain[307:304] ^ 1);
  assign w489[2] = |(datain[303:300] ^ 5);
  assign w489[3] = |(datain[299:296] ^ 6);
  assign w489[4] = |(datain[295:292] ^ 5);
  assign w489[5] = |(datain[291:288] ^ 7);
  assign w489[6] = |(datain[287:284] ^ 5);
  assign w489[7] = |(datain[283:280] ^ 3);
  assign w489[8] = |(datain[279:276] ^ 15);
  assign w489[9] = |(datain[275:272] ^ 15);
  assign w489[10] = |(datain[271:268] ^ 3);
  assign w489[11] = |(datain[267:264] ^ 6);
  assign w489[12] = |(datain[263:260] ^ 0);
  assign w489[13] = |(datain[259:256] ^ 12);
  assign w489[14] = |(datain[255:252] ^ 0);
  assign w489[15] = |(datain[251:248] ^ 1);
  assign w489[16] = |(datain[247:244] ^ 14);
  assign w489[17] = |(datain[243:240] ^ 11);
  assign w489[18] = |(datain[239:236] ^ 4);
  assign w489[19] = |(datain[235:232] ^ 12);
  assign comp[489] = ~(|w489);
  wire [44-1:0] w490;
  assign w490[0] = |(datain[311:308] ^ 0);
  assign w490[1] = |(datain[307:304] ^ 1);
  assign w490[2] = |(datain[303:300] ^ 9);
  assign w490[3] = |(datain[299:296] ^ 0);
  assign w490[4] = |(datain[295:292] ^ 8);
  assign w490[5] = |(datain[291:288] ^ 13);
  assign w490[6] = |(datain[287:284] ^ 9);
  assign w490[7] = |(datain[283:280] ^ 4);
  assign w490[8] = |(datain[279:276] ^ 0);
  assign w490[9] = |(datain[275:272] ^ 6);
  assign w490[10] = |(datain[271:268] ^ 0);
  assign w490[11] = |(datain[267:264] ^ 1);
  assign w490[12] = |(datain[263:260] ^ 11);
  assign w490[13] = |(datain[259:256] ^ 4);
  assign w490[14] = |(datain[255:252] ^ 4);
  assign w490[15] = |(datain[251:248] ^ 0);
  assign w490[16] = |(datain[247:244] ^ 12);
  assign w490[17] = |(datain[243:240] ^ 13);
  assign w490[18] = |(datain[239:236] ^ 2);
  assign w490[19] = |(datain[235:232] ^ 1);
  assign w490[20] = |(datain[231:228] ^ 7);
  assign w490[21] = |(datain[227:224] ^ 2);
  assign w490[22] = |(datain[223:220] ^ 2);
  assign w490[23] = |(datain[219:216] ^ 2);
  assign w490[24] = |(datain[215:212] ^ 5);
  assign w490[25] = |(datain[211:208] ^ 8);
  assign w490[26] = |(datain[207:204] ^ 0);
  assign w490[27] = |(datain[203:200] ^ 5);
  assign w490[28] = |(datain[199:196] ^ 4);
  assign w490[29] = |(datain[195:192] ^ 12);
  assign w490[30] = |(datain[191:188] ^ 0);
  assign w490[31] = |(datain[187:184] ^ 0);
  assign w490[32] = |(datain[183:180] ^ 12);
  assign w490[33] = |(datain[179:176] ^ 6);
  assign w490[34] = |(datain[175:172] ^ 0);
  assign w490[35] = |(datain[171:168] ^ 5);
  assign w490[36] = |(datain[167:164] ^ 14);
  assign w490[37] = |(datain[163:160] ^ 9);
  assign w490[38] = |(datain[159:156] ^ 8);
  assign w490[39] = |(datain[155:152] ^ 9);
  assign w490[40] = |(datain[151:148] ^ 4);
  assign w490[41] = |(datain[147:144] ^ 5);
  assign w490[42] = |(datain[143:140] ^ 0);
  assign w490[43] = |(datain[139:136] ^ 1);
  assign comp[490] = ~(|w490);
  wire [74-1:0] w491;
  assign w491[0] = |(datain[311:308] ^ 11);
  assign w491[1] = |(datain[307:304] ^ 4);
  assign w491[2] = |(datain[303:300] ^ 4);
  assign w491[3] = |(datain[299:296] ^ 0);
  assign w491[4] = |(datain[295:292] ^ 12);
  assign w491[5] = |(datain[291:288] ^ 13);
  assign w491[6] = |(datain[287:284] ^ 2);
  assign w491[7] = |(datain[283:280] ^ 1);
  assign w491[8] = |(datain[279:276] ^ 3);
  assign w491[9] = |(datain[275:272] ^ 2);
  assign w491[10] = |(datain[271:268] ^ 12);
  assign w491[11] = |(datain[267:264] ^ 0);
  assign w491[12] = |(datain[263:260] ^ 14);
  assign w491[13] = |(datain[259:256] ^ 8);
  assign w491[14] = |(datain[255:252] ^ 2);
  assign w491[15] = |(datain[251:248] ^ 14);
  assign w491[16] = |(datain[247:244] ^ 0);
  assign w491[17] = |(datain[243:240] ^ 0);
  assign w491[18] = |(datain[239:236] ^ 5);
  assign w491[19] = |(datain[235:232] ^ 8);
  assign w491[20] = |(datain[231:228] ^ 2);
  assign w491[21] = |(datain[227:224] ^ 13);
  assign w491[22] = |(datain[223:220] ^ 0);
  assign w491[23] = |(datain[219:216] ^ 3);
  assign w491[24] = |(datain[215:212] ^ 0);
  assign w491[25] = |(datain[211:208] ^ 0);
  assign w491[26] = |(datain[207:204] ^ 10);
  assign w491[27] = |(datain[203:200] ^ 3);
  assign w491[28] = |(datain[199:196] ^ 8);
  assign w491[29] = |(datain[195:192] ^ 14);
  assign w491[30] = |(datain[191:188] ^ 0);
  assign w491[31] = |(datain[187:184] ^ 0);
  assign w491[32] = |(datain[183:180] ^ 11);
  assign w491[33] = |(datain[179:176] ^ 9);
  assign w491[34] = |(datain[175:172] ^ 0);
  assign w491[35] = |(datain[171:168] ^ 3);
  assign w491[36] = |(datain[167:164] ^ 0);
  assign w491[37] = |(datain[163:160] ^ 0);
  assign w491[38] = |(datain[159:156] ^ 11);
  assign w491[39] = |(datain[155:152] ^ 10);
  assign w491[40] = |(datain[151:148] ^ 8);
  assign w491[41] = |(datain[147:144] ^ 13);
  assign w491[42] = |(datain[143:140] ^ 0);
  assign w491[43] = |(datain[139:136] ^ 0);
  assign w491[44] = |(datain[135:132] ^ 11);
  assign w491[45] = |(datain[131:128] ^ 4);
  assign w491[46] = |(datain[127:124] ^ 4);
  assign w491[47] = |(datain[123:120] ^ 0);
  assign w491[48] = |(datain[119:116] ^ 12);
  assign w491[49] = |(datain[115:112] ^ 13);
  assign w491[50] = |(datain[111:108] ^ 2);
  assign w491[51] = |(datain[107:104] ^ 1);
  assign w491[52] = |(datain[103:100] ^ 11);
  assign w491[53] = |(datain[99:96] ^ 0);
  assign w491[54] = |(datain[95:92] ^ 0);
  assign w491[55] = |(datain[91:88] ^ 2);
  assign w491[56] = |(datain[87:84] ^ 14);
  assign w491[57] = |(datain[83:80] ^ 8);
  assign w491[58] = |(datain[79:76] ^ 1);
  assign w491[59] = |(datain[75:72] ^ 8);
  assign w491[60] = |(datain[71:68] ^ 0);
  assign w491[61] = |(datain[67:64] ^ 0);
  assign w491[62] = |(datain[63:60] ^ 11);
  assign w491[63] = |(datain[59:56] ^ 9);
  assign w491[64] = |(datain[55:52] ^ 4);
  assign w491[65] = |(datain[51:48] ^ 7);
  assign w491[66] = |(datain[47:44] ^ 0);
  assign w491[67] = |(datain[43:40] ^ 2);
  assign w491[68] = |(datain[39:36] ^ 3);
  assign w491[69] = |(datain[35:32] ^ 3);
  assign w491[70] = |(datain[31:28] ^ 13);
  assign w491[71] = |(datain[27:24] ^ 2);
  assign w491[72] = |(datain[23:20] ^ 11);
  assign w491[73] = |(datain[19:16] ^ 4);
  assign comp[491] = ~(|w491);
  wire [76-1:0] w492;
  assign w492[0] = |(datain[311:308] ^ 12);
  assign w492[1] = |(datain[307:304] ^ 13);
  assign w492[2] = |(datain[303:300] ^ 2);
  assign w492[3] = |(datain[299:296] ^ 1);
  assign w492[4] = |(datain[295:292] ^ 3);
  assign w492[5] = |(datain[291:288] ^ 2);
  assign w492[6] = |(datain[287:284] ^ 12);
  assign w492[7] = |(datain[283:280] ^ 0);
  assign w492[8] = |(datain[279:276] ^ 14);
  assign w492[9] = |(datain[275:272] ^ 8);
  assign w492[10] = |(datain[271:268] ^ 2);
  assign w492[11] = |(datain[267:264] ^ 7);
  assign w492[12] = |(datain[263:260] ^ 0);
  assign w492[13] = |(datain[259:256] ^ 0);
  assign w492[14] = |(datain[255:252] ^ 5);
  assign w492[15] = |(datain[251:248] ^ 8);
  assign w492[16] = |(datain[247:244] ^ 2);
  assign w492[17] = |(datain[243:240] ^ 13);
  assign w492[18] = |(datain[239:236] ^ 0);
  assign w492[19] = |(datain[235:232] ^ 3);
  assign w492[20] = |(datain[231:228] ^ 0);
  assign w492[21] = |(datain[227:224] ^ 0);
  assign w492[22] = |(datain[223:220] ^ 10);
  assign w492[23] = |(datain[219:216] ^ 3);
  assign w492[24] = |(datain[215:212] ^ 8);
  assign w492[25] = |(datain[211:208] ^ 0);
  assign w492[26] = |(datain[207:204] ^ 0);
  assign w492[27] = |(datain[203:200] ^ 0);
  assign w492[28] = |(datain[199:196] ^ 11);
  assign w492[29] = |(datain[195:192] ^ 9);
  assign w492[30] = |(datain[191:188] ^ 0);
  assign w492[31] = |(datain[187:184] ^ 3);
  assign w492[32] = |(datain[183:180] ^ 0);
  assign w492[33] = |(datain[179:176] ^ 0);
  assign w492[34] = |(datain[175:172] ^ 11);
  assign w492[35] = |(datain[171:168] ^ 10);
  assign w492[36] = |(datain[167:164] ^ 7);
  assign w492[37] = |(datain[163:160] ^ 15);
  assign w492[38] = |(datain[159:156] ^ 0);
  assign w492[39] = |(datain[155:152] ^ 0);
  assign w492[40] = |(datain[151:148] ^ 11);
  assign w492[41] = |(datain[147:144] ^ 4);
  assign w492[42] = |(datain[143:140] ^ 4);
  assign w492[43] = |(datain[139:136] ^ 0);
  assign w492[44] = |(datain[135:132] ^ 12);
  assign w492[45] = |(datain[131:128] ^ 13);
  assign w492[46] = |(datain[127:124] ^ 2);
  assign w492[47] = |(datain[123:120] ^ 1);
  assign w492[48] = |(datain[119:116] ^ 11);
  assign w492[49] = |(datain[115:112] ^ 0);
  assign w492[50] = |(datain[111:108] ^ 0);
  assign w492[51] = |(datain[107:104] ^ 2);
  assign w492[52] = |(datain[103:100] ^ 14);
  assign w492[53] = |(datain[99:96] ^ 8);
  assign w492[54] = |(datain[95:92] ^ 1);
  assign w492[55] = |(datain[91:88] ^ 1);
  assign w492[56] = |(datain[87:84] ^ 0);
  assign w492[57] = |(datain[83:80] ^ 0);
  assign w492[58] = |(datain[79:76] ^ 11);
  assign w492[59] = |(datain[75:72] ^ 9);
  assign w492[60] = |(datain[71:68] ^ 8);
  assign w492[61] = |(datain[67:64] ^ 13);
  assign w492[62] = |(datain[63:60] ^ 0);
  assign w492[63] = |(datain[59:56] ^ 2);
  assign w492[64] = |(datain[55:52] ^ 3);
  assign w492[65] = |(datain[51:48] ^ 3);
  assign w492[66] = |(datain[47:44] ^ 13);
  assign w492[67] = |(datain[43:40] ^ 2);
  assign w492[68] = |(datain[39:36] ^ 11);
  assign w492[69] = |(datain[35:32] ^ 4);
  assign w492[70] = |(datain[31:28] ^ 4);
  assign w492[71] = |(datain[27:24] ^ 0);
  assign w492[72] = |(datain[23:20] ^ 12);
  assign w492[73] = |(datain[19:16] ^ 13);
  assign w492[74] = |(datain[15:12] ^ 2);
  assign w492[75] = |(datain[11:8] ^ 1);
  assign comp[492] = ~(|w492);
  wire [28-1:0] w493;
  assign w493[0] = |(datain[311:308] ^ 13);
  assign w493[1] = |(datain[307:304] ^ 1);
  assign w493[2] = |(datain[303:300] ^ 14);
  assign w493[3] = |(datain[299:296] ^ 0);
  assign w493[4] = |(datain[295:292] ^ 8);
  assign w493[5] = |(datain[291:288] ^ 0);
  assign w493[6] = |(datain[287:284] ^ 14);
  assign w493[7] = |(datain[283:280] ^ 4);
  assign w493[8] = |(datain[279:276] ^ 0);
  assign w493[9] = |(datain[275:272] ^ 3);
  assign w493[10] = |(datain[271:268] ^ 8);
  assign w493[11] = |(datain[267:264] ^ 0);
  assign w493[12] = |(datain[263:260] ^ 12);
  assign w493[13] = |(datain[259:256] ^ 4);
  assign w493[14] = |(datain[255:252] ^ 0);
  assign w493[15] = |(datain[251:248] ^ 2);
  assign w493[16] = |(datain[247:244] ^ 8);
  assign w493[17] = |(datain[243:240] ^ 10);
  assign w493[18] = |(datain[239:236] ^ 12);
  assign w493[19] = |(datain[235:232] ^ 4);
  assign w493[20] = |(datain[231:228] ^ 8);
  assign w493[21] = |(datain[227:224] ^ 11);
  assign w493[22] = |(datain[223:220] ^ 13);
  assign w493[23] = |(datain[219:216] ^ 8);
  assign w493[24] = |(datain[215:212] ^ 3);
  assign w493[25] = |(datain[211:208] ^ 2);
  assign w493[26] = |(datain[207:204] ^ 15);
  assign w493[27] = |(datain[203:200] ^ 15);
  assign comp[493] = ~(|w493);
  wire [30-1:0] w494;
  assign w494[0] = |(datain[311:308] ^ 11);
  assign w494[1] = |(datain[307:304] ^ 14);
  assign w494[2] = |(datain[303:300] ^ 0);
  assign w494[3] = |(datain[299:296] ^ 0);
  assign w494[4] = |(datain[295:292] ^ 0);
  assign w494[5] = |(datain[291:288] ^ 1);
  assign w494[6] = |(datain[287:284] ^ 5);
  assign w494[7] = |(datain[283:280] ^ 10);
  assign w494[8] = |(datain[279:276] ^ 5);
  assign w494[9] = |(datain[275:272] ^ 8);
  assign w494[10] = |(datain[271:268] ^ 15);
  assign w494[11] = |(datain[267:264] ^ 15);
  assign w494[12] = |(datain[263:260] ^ 14);
  assign w494[13] = |(datain[259:256] ^ 6);
  assign w494[14] = |(datain[255:252] ^ 5);
  assign w494[15] = |(datain[251:248] ^ 0);
  assign w494[16] = |(datain[247:244] ^ 11);
  assign w494[17] = |(datain[243:240] ^ 4);
  assign w494[18] = |(datain[239:236] ^ 0);
  assign w494[19] = |(datain[235:232] ^ 14);
  assign w494[20] = |(datain[231:228] ^ 8);
  assign w494[21] = |(datain[227:224] ^ 10);
  assign w494[22] = |(datain[223:220] ^ 13);
  assign w494[23] = |(datain[219:216] ^ 0);
  assign w494[24] = |(datain[215:212] ^ 12);
  assign w494[25] = |(datain[211:208] ^ 13);
  assign w494[26] = |(datain[207:204] ^ 2);
  assign w494[27] = |(datain[203:200] ^ 1);
  assign w494[28] = |(datain[199:196] ^ 5);
  assign w494[29] = |(datain[195:192] ^ 8);
  assign comp[494] = ~(|w494);
  wire [24-1:0] w495;
  assign w495[0] = |(datain[311:308] ^ 11);
  assign w495[1] = |(datain[307:304] ^ 0);
  assign w495[2] = |(datain[303:300] ^ 0);
  assign w495[3] = |(datain[299:296] ^ 0);
  assign w495[4] = |(datain[295:292] ^ 14);
  assign w495[5] = |(datain[291:288] ^ 8);
  assign w495[6] = |(datain[287:284] ^ 12);
  assign w495[7] = |(datain[283:280] ^ 0);
  assign w495[8] = |(datain[279:276] ^ 15);
  assign w495[9] = |(datain[275:272] ^ 15);
  assign w495[10] = |(datain[271:268] ^ 11);
  assign w495[11] = |(datain[267:264] ^ 4);
  assign w495[12] = |(datain[263:260] ^ 4);
  assign w495[13] = |(datain[259:256] ^ 0);
  assign w495[14] = |(datain[255:252] ^ 11);
  assign w495[15] = |(datain[251:248] ^ 10);
  assign w495[16] = |(datain[247:244] ^ 0);
  assign w495[17] = |(datain[243:240] ^ 0);
  assign w495[18] = |(datain[239:236] ^ 0);
  assign w495[19] = |(datain[235:232] ^ 1);
  assign w495[20] = |(datain[231:228] ^ 8);
  assign w495[21] = |(datain[227:224] ^ 11);
  assign w495[22] = |(datain[223:220] ^ 0);
  assign w495[23] = |(datain[219:216] ^ 14);
  assign comp[495] = ~(|w495);
  wire [42-1:0] w496;
  assign w496[0] = |(datain[311:308] ^ 14);
  assign w496[1] = |(datain[307:304] ^ 11);
  assign w496[2] = |(datain[303:300] ^ 1);
  assign w496[3] = |(datain[299:296] ^ 4);
  assign w496[4] = |(datain[295:292] ^ 11);
  assign w496[5] = |(datain[291:288] ^ 14);
  assign w496[6] = |(datain[287:284] ^ 3);
  assign w496[7] = |(datain[283:280] ^ 0);
  assign w496[8] = |(datain[279:276] ^ 0);
  assign w496[9] = |(datain[275:272] ^ 0);
  assign w496[10] = |(datain[271:268] ^ 0);
  assign w496[11] = |(datain[267:264] ^ 3);
  assign w496[12] = |(datain[263:260] ^ 15);
  assign w496[13] = |(datain[259:256] ^ 2);
  assign w496[14] = |(datain[255:252] ^ 8);
  assign w496[15] = |(datain[251:248] ^ 11);
  assign w496[16] = |(datain[247:244] ^ 15);
  assign w496[17] = |(datain[243:240] ^ 14);
  assign w496[18] = |(datain[239:236] ^ 8);
  assign w496[19] = |(datain[235:232] ^ 1);
  assign w496[20] = |(datain[231:228] ^ 14);
  assign w496[21] = |(datain[227:224] ^ 15);
  assign w496[22] = |(datain[223:220] ^ 4);
  assign w496[23] = |(datain[219:216] ^ 0);
  assign w496[24] = |(datain[215:212] ^ 0);
  assign w496[25] = |(datain[211:208] ^ 1);
  assign w496[26] = |(datain[207:204] ^ 11);
  assign w496[27] = |(datain[203:200] ^ 9);
  assign w496[28] = |(datain[199:196] ^ 11);
  assign w496[29] = |(datain[195:192] ^ 15);
  assign w496[30] = |(datain[191:188] ^ 0);
  assign w496[31] = |(datain[187:184] ^ 3);
  assign w496[32] = |(datain[183:180] ^ 3);
  assign w496[33] = |(datain[179:176] ^ 1);
  assign w496[34] = |(datain[175:172] ^ 3);
  assign w496[35] = |(datain[171:168] ^ 12);
  assign w496[36] = |(datain[167:164] ^ 4);
  assign w496[37] = |(datain[163:160] ^ 6);
  assign w496[38] = |(datain[159:156] ^ 14);
  assign w496[39] = |(datain[155:152] ^ 2);
  assign w496[40] = |(datain[151:148] ^ 15);
  assign w496[41] = |(datain[147:144] ^ 11);
  assign comp[496] = ~(|w496);
  wire [32-1:0] w497;
  assign w497[0] = |(datain[311:308] ^ 10);
  assign w497[1] = |(datain[307:304] ^ 1);
  assign w497[2] = |(datain[303:300] ^ 1);
  assign w497[3] = |(datain[299:296] ^ 3);
  assign w497[4] = |(datain[295:292] ^ 0);
  assign w497[5] = |(datain[291:288] ^ 4);
  assign w497[6] = |(datain[287:284] ^ 4);
  assign w497[7] = |(datain[283:280] ^ 8);
  assign w497[8] = |(datain[279:276] ^ 10);
  assign w497[9] = |(datain[275:272] ^ 3);
  assign w497[10] = |(datain[271:268] ^ 1);
  assign w497[11] = |(datain[267:264] ^ 3);
  assign w497[12] = |(datain[263:260] ^ 0);
  assign w497[13] = |(datain[259:256] ^ 4);
  assign w497[14] = |(datain[255:252] ^ 11);
  assign w497[15] = |(datain[251:248] ^ 1);
  assign w497[16] = |(datain[247:244] ^ 0);
  assign w497[17] = |(datain[243:240] ^ 6);
  assign w497[18] = |(datain[239:236] ^ 13);
  assign w497[19] = |(datain[235:232] ^ 3);
  assign w497[20] = |(datain[231:228] ^ 14);
  assign w497[21] = |(datain[227:224] ^ 0);
  assign w497[22] = |(datain[223:220] ^ 8);
  assign w497[23] = |(datain[219:216] ^ 14);
  assign w497[24] = |(datain[215:212] ^ 12);
  assign w497[25] = |(datain[211:208] ^ 0);
  assign w497[26] = |(datain[207:204] ^ 11);
  assign w497[27] = |(datain[203:200] ^ 9);
  assign w497[28] = |(datain[199:196] ^ 0);
  assign w497[29] = |(datain[195:192] ^ 0);
  assign w497[30] = |(datain[191:188] ^ 0);
  assign w497[31] = |(datain[187:184] ^ 2);
  assign comp[497] = ~(|w497);
  wire [76-1:0] w498;
  assign w498[0] = |(datain[311:308] ^ 12);
  assign w498[1] = |(datain[307:304] ^ 13);
  assign w498[2] = |(datain[303:300] ^ 2);
  assign w498[3] = |(datain[299:296] ^ 1);
  assign w498[4] = |(datain[295:292] ^ 11);
  assign w498[5] = |(datain[291:288] ^ 4);
  assign w498[6] = |(datain[287:284] ^ 4);
  assign w498[7] = |(datain[283:280] ^ 0);
  assign w498[8] = |(datain[279:276] ^ 11);
  assign w498[9] = |(datain[275:272] ^ 9);
  assign w498[10] = |(datain[271:268] ^ 1);
  assign w498[11] = |(datain[267:264] ^ 12);
  assign w498[12] = |(datain[263:260] ^ 0);
  assign w498[13] = |(datain[259:256] ^ 0);
  assign w498[14] = |(datain[255:252] ^ 0);
  assign w498[15] = |(datain[251:248] ^ 14);
  assign w498[16] = |(datain[247:244] ^ 1);
  assign w498[17] = |(datain[243:240] ^ 15);
  assign w498[18] = |(datain[239:236] ^ 11);
  assign w498[19] = |(datain[235:232] ^ 10);
  assign w498[20] = |(datain[231:228] ^ 4);
  assign w498[21] = |(datain[227:224] ^ 12);
  assign w498[22] = |(datain[223:220] ^ 0);
  assign w498[23] = |(datain[219:216] ^ 2);
  assign w498[24] = |(datain[215:212] ^ 12);
  assign w498[25] = |(datain[211:208] ^ 13);
  assign w498[26] = |(datain[207:204] ^ 2);
  assign w498[27] = |(datain[203:200] ^ 1);
  assign w498[28] = |(datain[199:196] ^ 5);
  assign w498[29] = |(datain[195:192] ^ 3);
  assign w498[30] = |(datain[191:188] ^ 6);
  assign w498[31] = |(datain[187:184] ^ 1);
  assign w498[32] = |(datain[183:180] ^ 6);
  assign w498[33] = |(datain[179:176] ^ 0);
  assign w498[34] = |(datain[175:172] ^ 5);
  assign w498[35] = |(datain[171:168] ^ 11);
  assign w498[36] = |(datain[167:164] ^ 6);
  assign w498[37] = |(datain[163:160] ^ 8);
  assign w498[38] = |(datain[159:156] ^ 0);
  assign w498[39] = |(datain[155:152] ^ 1);
  assign w498[40] = |(datain[151:148] ^ 5);
  assign w498[41] = |(datain[147:144] ^ 7);
  assign w498[42] = |(datain[143:140] ^ 5);
  assign w498[43] = |(datain[139:136] ^ 8);
  assign w498[44] = |(datain[135:132] ^ 2);
  assign w498[45] = |(datain[131:128] ^ 14);
  assign w498[46] = |(datain[127:124] ^ 8);
  assign w498[47] = |(datain[123:120] ^ 11);
  assign w498[48] = |(datain[119:116] ^ 0);
  assign w498[49] = |(datain[115:112] ^ 14);
  assign w498[50] = |(datain[111:108] ^ 4);
  assign w498[51] = |(datain[107:104] ^ 6);
  assign w498[52] = |(datain[103:100] ^ 0);
  assign w498[53] = |(datain[99:96] ^ 2);
  assign w498[54] = |(datain[95:92] ^ 2);
  assign w498[55] = |(datain[91:88] ^ 14);
  assign w498[56] = |(datain[87:84] ^ 8);
  assign w498[57] = |(datain[83:80] ^ 11);
  assign w498[58] = |(datain[79:76] ^ 1);
  assign w498[59] = |(datain[75:72] ^ 6);
  assign w498[60] = |(datain[71:68] ^ 4);
  assign w498[61] = |(datain[67:64] ^ 8);
  assign w498[62] = |(datain[63:60] ^ 0);
  assign w498[63] = |(datain[59:56] ^ 2);
  assign w498[64] = |(datain[55:52] ^ 12);
  assign w498[65] = |(datain[51:48] ^ 13);
  assign w498[66] = |(datain[47:44] ^ 2);
  assign w498[67] = |(datain[43:40] ^ 1);
  assign w498[68] = |(datain[39:36] ^ 11);
  assign w498[69] = |(datain[35:32] ^ 4);
  assign w498[70] = |(datain[31:28] ^ 3);
  assign w498[71] = |(datain[27:24] ^ 14);
  assign w498[72] = |(datain[23:20] ^ 12);
  assign w498[73] = |(datain[19:16] ^ 13);
  assign w498[74] = |(datain[15:12] ^ 2);
  assign w498[75] = |(datain[11:8] ^ 1);
  assign comp[498] = ~(|w498);
  wire [42-1:0] w499;
  assign w499[0] = |(datain[311:308] ^ 8);
  assign w499[1] = |(datain[307:304] ^ 14);
  assign w499[2] = |(datain[303:300] ^ 13);
  assign w499[3] = |(datain[299:296] ^ 8);
  assign w499[4] = |(datain[295:292] ^ 8);
  assign w499[5] = |(datain[291:288] ^ 0);
  assign w499[6] = |(datain[287:284] ^ 3);
  assign w499[7] = |(datain[283:280] ^ 14);
  assign w499[8] = |(datain[279:276] ^ 7);
  assign w499[9] = |(datain[275:272] ^ 2);
  assign w499[10] = |(datain[271:268] ^ 0);
  assign w499[11] = |(datain[267:264] ^ 4);
  assign w499[12] = |(datain[263:260] ^ 3);
  assign w499[13] = |(datain[259:256] ^ 12);
  assign w499[14] = |(datain[255:252] ^ 7);
  assign w499[15] = |(datain[251:248] ^ 4);
  assign w499[16] = |(datain[247:244] ^ 4);
  assign w499[17] = |(datain[243:240] ^ 8);
  assign w499[18] = |(datain[239:236] ^ 15);
  assign w499[19] = |(datain[235:232] ^ 10);
  assign w499[20] = |(datain[231:228] ^ 11);
  assign w499[21] = |(datain[227:224] ^ 14);
  assign w499[22] = |(datain[223:220] ^ 0);
  assign w499[23] = |(datain[219:216] ^ 3);
  assign w499[24] = |(datain[215:212] ^ 0);
  assign w499[25] = |(datain[211:208] ^ 4);
  assign w499[26] = |(datain[207:204] ^ 10);
  assign w499[27] = |(datain[203:200] ^ 13);
  assign w499[28] = |(datain[199:196] ^ 4);
  assign w499[29] = |(datain[195:192] ^ 8);
  assign w499[30] = |(datain[191:188] ^ 4);
  assign w499[31] = |(datain[187:184] ^ 14);
  assign w499[32] = |(datain[183:180] ^ 4);
  assign w499[33] = |(datain[179:176] ^ 14);
  assign w499[34] = |(datain[175:172] ^ 8);
  assign w499[35] = |(datain[171:168] ^ 9);
  assign w499[36] = |(datain[167:164] ^ 0);
  assign w499[37] = |(datain[163:160] ^ 4);
  assign w499[38] = |(datain[159:156] ^ 15);
  assign w499[39] = |(datain[155:152] ^ 11);
  assign w499[40] = |(datain[151:148] ^ 11);
  assign w499[41] = |(datain[147:144] ^ 1);
  assign comp[499] = ~(|w499);
  wire [46-1:0] w500;
  assign w500[0] = |(datain[311:308] ^ 8);
  assign w500[1] = |(datain[307:304] ^ 9);
  assign w500[2] = |(datain[303:300] ^ 8);
  assign w500[3] = |(datain[299:296] ^ 4);
  assign w500[4] = |(datain[295:292] ^ 1);
  assign w500[5] = |(datain[291:288] ^ 4);
  assign w500[6] = |(datain[287:284] ^ 0);
  assign w500[7] = |(datain[283:280] ^ 8);
  assign w500[8] = |(datain[279:276] ^ 11);
  assign w500[9] = |(datain[275:272] ^ 8);
  assign w500[10] = |(datain[271:268] ^ 0);
  assign w500[11] = |(datain[267:264] ^ 10);
  assign w500[12] = |(datain[263:260] ^ 0);
  assign w500[13] = |(datain[259:256] ^ 8);
  assign w500[14] = |(datain[255:252] ^ 0);
  assign w500[15] = |(datain[251:248] ^ 3);
  assign w500[16] = |(datain[247:244] ^ 12);
  assign w500[17] = |(datain[243:240] ^ 6);
  assign w500[18] = |(datain[239:236] ^ 10);
  assign w500[19] = |(datain[235:232] ^ 3);
  assign w500[20] = |(datain[231:228] ^ 0);
  assign w500[21] = |(datain[227:224] ^ 4);
  assign w500[22] = |(datain[223:220] ^ 0);
  assign w500[23] = |(datain[219:216] ^ 0);
  assign w500[24] = |(datain[215:212] ^ 8);
  assign w500[25] = |(datain[211:208] ^ 12);
  assign w500[26] = |(datain[207:204] ^ 0);
  assign w500[27] = |(datain[203:200] ^ 14);
  assign w500[28] = |(datain[199:196] ^ 0);
  assign w500[29] = |(datain[195:192] ^ 6);
  assign w500[30] = |(datain[191:188] ^ 0);
  assign w500[31] = |(datain[187:184] ^ 0);
  assign w500[32] = |(datain[183:180] ^ 9);
  assign w500[33] = |(datain[179:176] ^ 12);
  assign w500[34] = |(datain[175:172] ^ 5);
  assign w500[35] = |(datain[171:168] ^ 8);
  assign w500[36] = |(datain[167:164] ^ 0);
  assign w500[37] = |(datain[163:160] ^ 13);
  assign w500[38] = |(datain[159:156] ^ 0);
  assign w500[39] = |(datain[155:152] ^ 0);
  assign w500[40] = |(datain[151:148] ^ 0);
  assign w500[41] = |(datain[147:144] ^ 1);
  assign w500[42] = |(datain[143:140] ^ 5);
  assign w500[43] = |(datain[139:136] ^ 0);
  assign w500[44] = |(datain[135:132] ^ 9);
  assign w500[45] = |(datain[131:128] ^ 13);
  assign comp[500] = ~(|w500);
  wire [40-1:0] w501;
  assign w501[0] = |(datain[311:308] ^ 8);
  assign w501[1] = |(datain[307:304] ^ 7);
  assign w501[2] = |(datain[303:300] ^ 12);
  assign w501[3] = |(datain[299:296] ^ 15);
  assign w501[4] = |(datain[295:292] ^ 12);
  assign w501[5] = |(datain[291:288] ^ 13);
  assign w501[6] = |(datain[287:284] ^ 2);
  assign w501[7] = |(datain[283:280] ^ 1);
  assign w501[8] = |(datain[279:276] ^ 11);
  assign w501[9] = |(datain[275:272] ^ 4);
  assign w501[10] = |(datain[271:268] ^ 4);
  assign w501[11] = |(datain[267:264] ^ 0);
  assign w501[12] = |(datain[263:260] ^ 5);
  assign w501[13] = |(datain[259:256] ^ 10);
  assign w501[14] = |(datain[255:252] ^ 8);
  assign w501[15] = |(datain[251:248] ^ 7);
  assign w501[16] = |(datain[247:244] ^ 12);
  assign w501[17] = |(datain[243:240] ^ 15);
  assign w501[18] = |(datain[239:236] ^ 12);
  assign w501[19] = |(datain[235:232] ^ 13);
  assign w501[20] = |(datain[231:228] ^ 2);
  assign w501[21] = |(datain[227:224] ^ 1);
  assign w501[22] = |(datain[223:220] ^ 11);
  assign w501[23] = |(datain[219:216] ^ 4);
  assign w501[24] = |(datain[215:212] ^ 3);
  assign w501[25] = |(datain[211:208] ^ 14);
  assign w501[26] = |(datain[207:204] ^ 12);
  assign w501[27] = |(datain[203:200] ^ 13);
  assign w501[28] = |(datain[199:196] ^ 2);
  assign w501[29] = |(datain[195:192] ^ 1);
  assign w501[30] = |(datain[191:188] ^ 11);
  assign w501[31] = |(datain[187:184] ^ 4);
  assign w501[32] = |(datain[183:180] ^ 4);
  assign w501[33] = |(datain[179:176] ^ 15);
  assign w501[34] = |(datain[175:172] ^ 12);
  assign w501[35] = |(datain[171:168] ^ 13);
  assign w501[36] = |(datain[167:164] ^ 2);
  assign w501[37] = |(datain[163:160] ^ 1);
  assign w501[38] = |(datain[159:156] ^ 7);
  assign w501[39] = |(datain[155:152] ^ 3);
  assign comp[501] = ~(|w501);
  wire [28-1:0] w502;
  assign w502[0] = |(datain[311:308] ^ 11);
  assign w502[1] = |(datain[307:304] ^ 10);
  assign w502[2] = |(datain[303:300] ^ 15);
  assign w502[3] = |(datain[299:296] ^ 2);
  assign w502[4] = |(datain[295:292] ^ 0);
  assign w502[5] = |(datain[291:288] ^ 0);
  assign w502[6] = |(datain[287:284] ^ 11);
  assign w502[7] = |(datain[283:280] ^ 8);
  assign w502[8] = |(datain[279:276] ^ 0);
  assign w502[9] = |(datain[275:272] ^ 2);
  assign w502[10] = |(datain[271:268] ^ 3);
  assign w502[11] = |(datain[267:264] ^ 13);
  assign w502[12] = |(datain[263:260] ^ 12);
  assign w502[13] = |(datain[259:256] ^ 13);
  assign w502[14] = |(datain[255:252] ^ 2);
  assign w502[15] = |(datain[251:248] ^ 1);
  assign w502[16] = |(datain[247:244] ^ 8);
  assign w502[17] = |(datain[243:240] ^ 11);
  assign w502[18] = |(datain[239:236] ^ 13);
  assign w502[19] = |(datain[235:232] ^ 8);
  assign w502[20] = |(datain[231:228] ^ 7);
  assign w502[21] = |(datain[227:224] ^ 2);
  assign w502[22] = |(datain[223:220] ^ 3);
  assign w502[23] = |(datain[219:216] ^ 4);
  assign w502[24] = |(datain[215:212] ^ 11);
  assign w502[25] = |(datain[211:208] ^ 4);
  assign w502[26] = |(datain[207:204] ^ 3);
  assign w502[27] = |(datain[203:200] ^ 15);
  assign comp[502] = ~(|w502);
  wire [48-1:0] w503;
  assign w503[0] = |(datain[311:308] ^ 11);
  assign w503[1] = |(datain[307:304] ^ 8);
  assign w503[2] = |(datain[303:300] ^ 0);
  assign w503[3] = |(datain[299:296] ^ 0);
  assign w503[4] = |(datain[295:292] ^ 4);
  assign w503[5] = |(datain[291:288] ^ 2);
  assign w503[6] = |(datain[287:284] ^ 5);
  assign w503[7] = |(datain[283:280] ^ 10);
  assign w503[8] = |(datain[279:276] ^ 8);
  assign w503[9] = |(datain[275:272] ^ 7);
  assign w503[10] = |(datain[271:268] ^ 12);
  assign w503[11] = |(datain[267:264] ^ 15);
  assign w503[12] = |(datain[263:260] ^ 12);
  assign w503[13] = |(datain[259:256] ^ 13);
  assign w503[14] = |(datain[255:252] ^ 2);
  assign w503[15] = |(datain[251:248] ^ 1);
  assign w503[16] = |(datain[247:244] ^ 11);
  assign w503[17] = |(datain[243:240] ^ 4);
  assign w503[18] = |(datain[239:236] ^ 4);
  assign w503[19] = |(datain[235:232] ^ 0);
  assign w503[20] = |(datain[231:228] ^ 5);
  assign w503[21] = |(datain[227:224] ^ 10);
  assign w503[22] = |(datain[223:220] ^ 8);
  assign w503[23] = |(datain[219:216] ^ 7);
  assign w503[24] = |(datain[215:212] ^ 12);
  assign w503[25] = |(datain[211:208] ^ 15);
  assign w503[26] = |(datain[207:204] ^ 12);
  assign w503[27] = |(datain[203:200] ^ 13);
  assign w503[28] = |(datain[199:196] ^ 2);
  assign w503[29] = |(datain[195:192] ^ 1);
  assign w503[30] = |(datain[191:188] ^ 11);
  assign w503[31] = |(datain[187:184] ^ 4);
  assign w503[32] = |(datain[183:180] ^ 3);
  assign w503[33] = |(datain[179:176] ^ 14);
  assign w503[34] = |(datain[175:172] ^ 12);
  assign w503[35] = |(datain[171:168] ^ 13);
  assign w503[36] = |(datain[167:164] ^ 2);
  assign w503[37] = |(datain[163:160] ^ 1);
  assign w503[38] = |(datain[159:156] ^ 11);
  assign w503[39] = |(datain[155:152] ^ 4);
  assign w503[40] = |(datain[151:148] ^ 4);
  assign w503[41] = |(datain[147:144] ^ 15);
  assign w503[42] = |(datain[143:140] ^ 12);
  assign w503[43] = |(datain[139:136] ^ 13);
  assign w503[44] = |(datain[135:132] ^ 2);
  assign w503[45] = |(datain[131:128] ^ 1);
  assign w503[46] = |(datain[127:124] ^ 7);
  assign w503[47] = |(datain[123:120] ^ 3);
  assign comp[503] = ~(|w503);
  wire [76-1:0] w504;
  assign w504[0] = |(datain[311:308] ^ 0);
  assign w504[1] = |(datain[307:304] ^ 1);
  assign w504[2] = |(datain[303:300] ^ 7);
  assign w504[3] = |(datain[299:296] ^ 2);
  assign w504[4] = |(datain[295:292] ^ 2);
  assign w504[5] = |(datain[291:288] ^ 14);
  assign w504[6] = |(datain[287:284] ^ 3);
  assign w504[7] = |(datain[283:280] ^ 13);
  assign w504[8] = |(datain[279:276] ^ 7);
  assign w504[9] = |(datain[275:272] ^ 0);
  assign w504[10] = |(datain[271:268] ^ 15);
  assign w504[11] = |(datain[267:264] ^ 11);
  assign w504[12] = |(datain[263:260] ^ 7);
  assign w504[13] = |(datain[259:256] ^ 7);
  assign w504[14] = |(datain[255:252] ^ 2);
  assign w504[15] = |(datain[251:248] ^ 9);
  assign w504[16] = |(datain[247:244] ^ 2);
  assign w504[17] = |(datain[243:240] ^ 13);
  assign w504[18] = |(datain[239:236] ^ 0);
  assign w504[19] = |(datain[235:232] ^ 3);
  assign w504[20] = |(datain[231:228] ^ 0);
  assign w504[21] = |(datain[227:224] ^ 0);
  assign w504[22] = |(datain[223:220] ^ 2);
  assign w504[23] = |(datain[219:216] ^ 14);
  assign w504[24] = |(datain[215:212] ^ 10);
  assign w504[25] = |(datain[211:208] ^ 3);
  assign w504[26] = |(datain[207:204] ^ 0);
  assign w504[27] = |(datain[203:200] ^ 14);
  assign w504[28] = |(datain[199:196] ^ 0);
  assign w504[29] = |(datain[195:192] ^ 1);
  assign w504[30] = |(datain[191:188] ^ 11);
  assign w504[31] = |(datain[187:184] ^ 4);
  assign w504[32] = |(datain[183:180] ^ 4);
  assign w504[33] = |(datain[179:176] ^ 0);
  assign w504[34] = |(datain[175:172] ^ 11);
  assign w504[35] = |(datain[171:168] ^ 9);
  assign w504[36] = |(datain[167:164] ^ 1);
  assign w504[37] = |(datain[163:160] ^ 0);
  assign w504[38] = |(datain[159:156] ^ 0);
  assign w504[39] = |(datain[155:152] ^ 3);
  assign w504[40] = |(datain[151:148] ^ 9);
  assign w504[41] = |(datain[147:144] ^ 0);
  assign w504[42] = |(datain[143:140] ^ 11);
  assign w504[43] = |(datain[139:136] ^ 10);
  assign w504[44] = |(datain[135:132] ^ 0);
  assign w504[45] = |(datain[131:128] ^ 0);
  assign w504[46] = |(datain[127:124] ^ 0);
  assign w504[47] = |(datain[123:120] ^ 1);
  assign w504[48] = |(datain[119:116] ^ 12);
  assign w504[49] = |(datain[115:112] ^ 13);
  assign w504[50] = |(datain[111:108] ^ 2);
  assign w504[51] = |(datain[107:104] ^ 1);
  assign w504[52] = |(datain[103:100] ^ 7);
  assign w504[53] = |(datain[99:96] ^ 2);
  assign w504[54] = |(datain[95:92] ^ 1);
  assign w504[55] = |(datain[91:88] ^ 5);
  assign w504[56] = |(datain[87:84] ^ 11);
  assign w504[57] = |(datain[83:80] ^ 8);
  assign w504[58] = |(datain[79:76] ^ 0);
  assign w504[59] = |(datain[75:72] ^ 0);
  assign w504[60] = |(datain[71:68] ^ 4);
  assign w504[61] = |(datain[67:64] ^ 2);
  assign w504[62] = |(datain[63:60] ^ 3);
  assign w504[63] = |(datain[59:56] ^ 3);
  assign w504[64] = |(datain[55:52] ^ 12);
  assign w504[65] = |(datain[51:48] ^ 9);
  assign w504[66] = |(datain[47:44] ^ 3);
  assign w504[67] = |(datain[43:40] ^ 3);
  assign w504[68] = |(datain[39:36] ^ 13);
  assign w504[69] = |(datain[35:32] ^ 2);
  assign w504[70] = |(datain[31:28] ^ 12);
  assign w504[71] = |(datain[27:24] ^ 13);
  assign w504[72] = |(datain[23:20] ^ 2);
  assign w504[73] = |(datain[19:16] ^ 1);
  assign w504[74] = |(datain[15:12] ^ 7);
  assign w504[75] = |(datain[11:8] ^ 2);
  assign comp[504] = ~(|w504);
  wire [64-1:0] w505;
  assign w505[0] = |(datain[311:308] ^ 8);
  assign w505[1] = |(datain[307:304] ^ 11);
  assign w505[2] = |(datain[303:300] ^ 8);
  assign w505[3] = |(datain[299:296] ^ 6);
  assign w505[4] = |(datain[295:292] ^ 8);
  assign w505[5] = |(datain[291:288] ^ 2);
  assign w505[6] = |(datain[287:284] ^ 0);
  assign w505[7] = |(datain[283:280] ^ 1);
  assign w505[8] = |(datain[279:276] ^ 3);
  assign w505[9] = |(datain[275:272] ^ 1);
  assign w505[10] = |(datain[271:268] ^ 0);
  assign w505[11] = |(datain[267:264] ^ 7);
  assign w505[12] = |(datain[263:260] ^ 4);
  assign w505[13] = |(datain[259:256] ^ 3);
  assign w505[14] = |(datain[255:252] ^ 4);
  assign w505[15] = |(datain[251:248] ^ 3);
  assign w505[16] = |(datain[247:244] ^ 14);
  assign w505[17] = |(datain[243:240] ^ 2);
  assign w505[18] = |(datain[239:236] ^ 15);
  assign w505[19] = |(datain[235:232] ^ 10);
  assign w505[20] = |(datain[231:228] ^ 5);
  assign w505[21] = |(datain[227:224] ^ 11);
  assign w505[22] = |(datain[223:220] ^ 12);
  assign w505[23] = |(datain[219:216] ^ 3);
  assign w505[24] = |(datain[215:212] ^ 14);
  assign w505[25] = |(datain[211:208] ^ 8);
  assign w505[26] = |(datain[207:204] ^ 14);
  assign w505[27] = |(datain[203:200] ^ 9);
  assign w505[28] = |(datain[199:196] ^ 15);
  assign w505[29] = |(datain[195:192] ^ 15);
  assign w505[30] = |(datain[191:188] ^ 11);
  assign w505[31] = |(datain[187:184] ^ 4);
  assign w505[32] = |(datain[183:180] ^ 4);
  assign w505[33] = |(datain[179:176] ^ 0);
  assign w505[34] = |(datain[175:172] ^ 8);
  assign w505[35] = |(datain[171:168] ^ 13);
  assign w505[36] = |(datain[167:164] ^ 9);
  assign w505[37] = |(datain[163:160] ^ 6);
  assign w505[38] = |(datain[159:156] ^ 0);
  assign w505[39] = |(datain[155:152] ^ 6);
  assign w505[40] = |(datain[151:148] ^ 0);
  assign w505[41] = |(datain[147:144] ^ 0);
  assign w505[42] = |(datain[143:140] ^ 11);
  assign w505[43] = |(datain[139:136] ^ 9);
  assign w505[44] = |(datain[135:132] ^ 8);
  assign w505[45] = |(datain[131:128] ^ 1);
  assign w505[46] = |(datain[127:124] ^ 0);
  assign w505[47] = |(datain[123:120] ^ 1);
  assign w505[48] = |(datain[119:116] ^ 12);
  assign w505[49] = |(datain[115:112] ^ 13);
  assign w505[50] = |(datain[111:108] ^ 2);
  assign w505[51] = |(datain[107:104] ^ 1);
  assign w505[52] = |(datain[103:100] ^ 14);
  assign w505[53] = |(datain[99:96] ^ 8);
  assign w505[54] = |(datain[95:92] ^ 13);
  assign w505[55] = |(datain[91:88] ^ 11);
  assign w505[56] = |(datain[87:84] ^ 15);
  assign w505[57] = |(datain[83:80] ^ 15);
  assign w505[58] = |(datain[79:76] ^ 12);
  assign w505[59] = |(datain[75:72] ^ 3);
  assign w505[60] = |(datain[71:68] ^ 7);
  assign w505[61] = |(datain[67:64] ^ 9);
  assign w505[62] = |(datain[63:60] ^ 6);
  assign w505[63] = |(datain[59:56] ^ 8);
  assign comp[505] = ~(|w505);
  wire [76-1:0] w506;
  assign w506[0] = |(datain[311:308] ^ 11);
  assign w506[1] = |(datain[307:304] ^ 9);
  assign w506[2] = |(datain[303:300] ^ 0);
  assign w506[3] = |(datain[299:296] ^ 2);
  assign w506[4] = |(datain[295:292] ^ 0);
  assign w506[5] = |(datain[291:288] ^ 0);
  assign w506[6] = |(datain[287:284] ^ 11);
  assign w506[7] = |(datain[283:280] ^ 10);
  assign w506[8] = |(datain[279:276] ^ 2);
  assign w506[9] = |(datain[275:272] ^ 9);
  assign w506[10] = |(datain[271:268] ^ 0);
  assign w506[11] = |(datain[267:264] ^ 1);
  assign w506[12] = |(datain[263:260] ^ 12);
  assign w506[13] = |(datain[259:256] ^ 13);
  assign w506[14] = |(datain[255:252] ^ 2);
  assign w506[15] = |(datain[251:248] ^ 1);
  assign w506[16] = |(datain[247:244] ^ 11);
  assign w506[17] = |(datain[243:240] ^ 8);
  assign w506[18] = |(datain[239:236] ^ 0);
  assign w506[19] = |(datain[235:232] ^ 2);
  assign w506[20] = |(datain[231:228] ^ 4);
  assign w506[21] = |(datain[227:224] ^ 2);
  assign w506[22] = |(datain[223:220] ^ 3);
  assign w506[23] = |(datain[219:216] ^ 3);
  assign w506[24] = |(datain[215:212] ^ 12);
  assign w506[25] = |(datain[211:208] ^ 9);
  assign w506[26] = |(datain[207:204] ^ 8);
  assign w506[27] = |(datain[203:200] ^ 11);
  assign w506[28] = |(datain[199:196] ^ 13);
  assign w506[29] = |(datain[195:192] ^ 1);
  assign w506[30] = |(datain[191:188] ^ 12);
  assign w506[31] = |(datain[187:184] ^ 13);
  assign w506[32] = |(datain[183:180] ^ 2);
  assign w506[33] = |(datain[179:176] ^ 1);
  assign w506[34] = |(datain[175:172] ^ 11);
  assign w506[35] = |(datain[171:168] ^ 9);
  assign w506[36] = |(datain[167:164] ^ 3);
  assign w506[37] = |(datain[163:160] ^ 6);
  assign w506[38] = |(datain[159:156] ^ 0);
  assign w506[39] = |(datain[155:152] ^ 8);
  assign w506[40] = |(datain[151:148] ^ 11);
  assign w506[41] = |(datain[147:144] ^ 4);
  assign w506[42] = |(datain[143:140] ^ 4);
  assign w506[43] = |(datain[139:136] ^ 0);
  assign w506[44] = |(datain[135:132] ^ 11);
  assign w506[45] = |(datain[131:128] ^ 10);
  assign w506[46] = |(datain[127:124] ^ 0);
  assign w506[47] = |(datain[123:120] ^ 0);
  assign w506[48] = |(datain[119:116] ^ 0);
  assign w506[49] = |(datain[115:112] ^ 1);
  assign w506[50] = |(datain[111:108] ^ 12);
  assign w506[51] = |(datain[107:104] ^ 13);
  assign w506[52] = |(datain[103:100] ^ 2);
  assign w506[53] = |(datain[99:96] ^ 1);
  assign w506[54] = |(datain[95:92] ^ 11);
  assign w506[55] = |(datain[91:88] ^ 10);
  assign w506[56] = |(datain[87:84] ^ 4);
  assign w506[57] = |(datain[83:80] ^ 8);
  assign w506[58] = |(datain[79:76] ^ 0);
  assign w506[59] = |(datain[75:72] ^ 1);
  assign w506[60] = |(datain[71:68] ^ 11);
  assign w506[61] = |(datain[67:64] ^ 9);
  assign w506[62] = |(datain[63:60] ^ 0);
  assign w506[63] = |(datain[59:56] ^ 6);
  assign w506[64] = |(datain[55:52] ^ 0);
  assign w506[65] = |(datain[51:48] ^ 0);
  assign w506[66] = |(datain[47:44] ^ 11);
  assign w506[67] = |(datain[43:40] ^ 4);
  assign w506[68] = |(datain[39:36] ^ 4);
  assign w506[69] = |(datain[35:32] ^ 0);
  assign w506[70] = |(datain[31:28] ^ 12);
  assign w506[71] = |(datain[27:24] ^ 13);
  assign w506[72] = |(datain[23:20] ^ 2);
  assign w506[73] = |(datain[19:16] ^ 1);
  assign w506[74] = |(datain[15:12] ^ 11);
  assign w506[75] = |(datain[11:8] ^ 8);
  assign comp[506] = ~(|w506);
  wire [46-1:0] w507;
  assign w507[0] = |(datain[311:308] ^ 5);
  assign w507[1] = |(datain[307:304] ^ 14);
  assign w507[2] = |(datain[303:300] ^ 13);
  assign w507[3] = |(datain[299:296] ^ 0);
  assign w507[4] = |(datain[295:292] ^ 12);
  assign w507[5] = |(datain[291:288] ^ 0);
  assign w507[6] = |(datain[287:284] ^ 11);
  assign w507[7] = |(datain[283:280] ^ 9);
  assign w507[8] = |(datain[279:276] ^ 3);
  assign w507[9] = |(datain[275:272] ^ 11);
  assign w507[10] = |(datain[271:268] ^ 0);
  assign w507[11] = |(datain[267:264] ^ 3);
  assign w507[12] = |(datain[263:260] ^ 15);
  assign w507[13] = |(datain[259:256] ^ 14);
  assign w507[14] = |(datain[255:252] ^ 12);
  assign w507[15] = |(datain[251:248] ^ 0);
  assign w507[16] = |(datain[247:244] ^ 2);
  assign w507[17] = |(datain[243:240] ^ 14);
  assign w507[18] = |(datain[239:236] ^ 8);
  assign w507[19] = |(datain[235:232] ^ 1);
  assign w507[20] = |(datain[231:228] ^ 3);
  assign w507[21] = |(datain[227:224] ^ 4);
  assign w507[22] = |(datain[223:220] ^ 1);
  assign w507[23] = |(datain[219:216] ^ 1);
  assign w507[24] = |(datain[215:212] ^ 9);
  assign w507[25] = |(datain[211:208] ^ 2);
  assign w507[26] = |(datain[207:204] ^ 15);
  assign w507[27] = |(datain[203:200] ^ 14);
  assign w507[28] = |(datain[199:196] ^ 12);
  assign w507[29] = |(datain[195:192] ^ 4);
  assign w507[30] = |(datain[191:188] ^ 4);
  assign w507[31] = |(datain[187:184] ^ 6);
  assign w507[32] = |(datain[183:180] ^ 15);
  assign w507[33] = |(datain[179:176] ^ 14);
  assign w507[34] = |(datain[175:172] ^ 12);
  assign w507[35] = |(datain[171:168] ^ 2);
  assign w507[36] = |(datain[167:164] ^ 4);
  assign w507[37] = |(datain[163:160] ^ 6);
  assign w507[38] = |(datain[159:156] ^ 13);
  assign w507[39] = |(datain[155:152] ^ 0);
  assign w507[40] = |(datain[151:148] ^ 12);
  assign w507[41] = |(datain[147:144] ^ 0);
  assign w507[42] = |(datain[143:140] ^ 14);
  assign w507[43] = |(datain[139:136] ^ 2);
  assign w507[44] = |(datain[135:132] ^ 15);
  assign w507[45] = |(datain[131:128] ^ 1);
  assign comp[507] = ~(|w507);
  wire [74-1:0] w508;
  assign w508[0] = |(datain[311:308] ^ 0);
  assign w508[1] = |(datain[307:304] ^ 3);
  assign w508[2] = |(datain[303:300] ^ 13);
  assign w508[3] = |(datain[299:296] ^ 6);
  assign w508[4] = |(datain[295:292] ^ 11);
  assign w508[5] = |(datain[291:288] ^ 9);
  assign w508[6] = |(datain[287:284] ^ 0);
  assign w508[7] = |(datain[283:280] ^ 14);
  assign w508[8] = |(datain[279:276] ^ 1);
  assign w508[9] = |(datain[275:272] ^ 1);
  assign w508[10] = |(datain[271:268] ^ 11);
  assign w508[11] = |(datain[267:264] ^ 4);
  assign w508[12] = |(datain[263:260] ^ 4);
  assign w508[13] = |(datain[259:256] ^ 0);
  assign w508[14] = |(datain[255:252] ^ 8);
  assign w508[15] = |(datain[251:248] ^ 11);
  assign w508[16] = |(datain[247:244] ^ 9);
  assign w508[17] = |(datain[243:240] ^ 12);
  assign w508[18] = |(datain[239:236] ^ 7);
  assign w508[19] = |(datain[235:232] ^ 4);
  assign w508[20] = |(datain[231:228] ^ 1);
  assign w508[21] = |(datain[227:224] ^ 2);
  assign w508[22] = |(datain[223:220] ^ 12);
  assign w508[23] = |(datain[219:216] ^ 13);
  assign w508[24] = |(datain[215:212] ^ 2);
  assign w508[25] = |(datain[211:208] ^ 1);
  assign w508[26] = |(datain[207:204] ^ 11);
  assign w508[27] = |(datain[203:200] ^ 8);
  assign w508[28] = |(datain[199:196] ^ 0);
  assign w508[29] = |(datain[195:192] ^ 0);
  assign w508[30] = |(datain[191:188] ^ 4);
  assign w508[31] = |(datain[187:184] ^ 2);
  assign w508[32] = |(datain[183:180] ^ 8);
  assign w508[33] = |(datain[179:176] ^ 11);
  assign w508[34] = |(datain[175:172] ^ 9);
  assign w508[35] = |(datain[171:168] ^ 12);
  assign w508[36] = |(datain[167:164] ^ 7);
  assign w508[37] = |(datain[163:160] ^ 4);
  assign w508[38] = |(datain[159:156] ^ 1);
  assign w508[39] = |(datain[155:152] ^ 2);
  assign w508[40] = |(datain[151:148] ^ 11);
  assign w508[41] = |(datain[147:144] ^ 9);
  assign w508[42] = |(datain[143:140] ^ 0);
  assign w508[43] = |(datain[139:136] ^ 0);
  assign w508[44] = |(datain[135:132] ^ 0);
  assign w508[45] = |(datain[131:128] ^ 0);
  assign w508[46] = |(datain[127:124] ^ 11);
  assign w508[47] = |(datain[123:120] ^ 10);
  assign w508[48] = |(datain[119:116] ^ 0);
  assign w508[49] = |(datain[115:112] ^ 0);
  assign w508[50] = |(datain[111:108] ^ 0);
  assign w508[51] = |(datain[107:104] ^ 0);
  assign w508[52] = |(datain[103:100] ^ 12);
  assign w508[53] = |(datain[99:96] ^ 13);
  assign w508[54] = |(datain[95:92] ^ 2);
  assign w508[55] = |(datain[91:88] ^ 1);
  assign w508[56] = |(datain[87:84] ^ 11);
  assign w508[57] = |(datain[83:80] ^ 4);
  assign w508[58] = |(datain[79:76] ^ 4);
  assign w508[59] = |(datain[75:72] ^ 0);
  assign w508[60] = |(datain[71:68] ^ 8);
  assign w508[61] = |(datain[67:64] ^ 11);
  assign w508[62] = |(datain[63:60] ^ 9);
  assign w508[63] = |(datain[59:56] ^ 12);
  assign w508[64] = |(datain[55:52] ^ 7);
  assign w508[65] = |(datain[51:48] ^ 4);
  assign w508[66] = |(datain[47:44] ^ 1);
  assign w508[67] = |(datain[43:40] ^ 2);
  assign w508[68] = |(datain[39:36] ^ 11);
  assign w508[69] = |(datain[35:32] ^ 9);
  assign w508[70] = |(datain[31:28] ^ 2);
  assign w508[71] = |(datain[27:24] ^ 0);
  assign w508[72] = |(datain[23:20] ^ 0);
  assign w508[73] = |(datain[19:16] ^ 0);
  assign comp[508] = ~(|w508);
  wire [72-1:0] w509;
  assign w509[0] = |(datain[311:308] ^ 13);
  assign w509[1] = |(datain[307:304] ^ 6);
  assign w509[2] = |(datain[303:300] ^ 11);
  assign w509[3] = |(datain[299:296] ^ 9);
  assign w509[4] = |(datain[295:292] ^ 11);
  assign w509[5] = |(datain[291:288] ^ 7);
  assign w509[6] = |(datain[287:284] ^ 0);
  assign w509[7] = |(datain[283:280] ^ 2);
  assign w509[8] = |(datain[279:276] ^ 11);
  assign w509[9] = |(datain[275:272] ^ 4);
  assign w509[10] = |(datain[271:268] ^ 4);
  assign w509[11] = |(datain[267:264] ^ 0);
  assign w509[12] = |(datain[263:260] ^ 8);
  assign w509[13] = |(datain[259:256] ^ 11);
  assign w509[14] = |(datain[255:252] ^ 9);
  assign w509[15] = |(datain[251:248] ^ 12);
  assign w509[16] = |(datain[247:244] ^ 6);
  assign w509[17] = |(datain[243:240] ^ 2);
  assign w509[18] = |(datain[239:236] ^ 0);
  assign w509[19] = |(datain[235:232] ^ 6);
  assign w509[20] = |(datain[231:228] ^ 12);
  assign w509[21] = |(datain[227:224] ^ 13);
  assign w509[22] = |(datain[223:220] ^ 2);
  assign w509[23] = |(datain[219:216] ^ 1);
  assign w509[24] = |(datain[215:212] ^ 11);
  assign w509[25] = |(datain[211:208] ^ 8);
  assign w509[26] = |(datain[207:204] ^ 0);
  assign w509[27] = |(datain[203:200] ^ 0);
  assign w509[28] = |(datain[199:196] ^ 4);
  assign w509[29] = |(datain[195:192] ^ 2);
  assign w509[30] = |(datain[191:188] ^ 8);
  assign w509[31] = |(datain[187:184] ^ 11);
  assign w509[32] = |(datain[183:180] ^ 9);
  assign w509[33] = |(datain[179:176] ^ 12);
  assign w509[34] = |(datain[175:172] ^ 6);
  assign w509[35] = |(datain[171:168] ^ 2);
  assign w509[36] = |(datain[167:164] ^ 0);
  assign w509[37] = |(datain[163:160] ^ 6);
  assign w509[38] = |(datain[159:156] ^ 11);
  assign w509[39] = |(datain[155:152] ^ 9);
  assign w509[40] = |(datain[151:148] ^ 0);
  assign w509[41] = |(datain[147:144] ^ 0);
  assign w509[42] = |(datain[143:140] ^ 0);
  assign w509[43] = |(datain[139:136] ^ 0);
  assign w509[44] = |(datain[135:132] ^ 11);
  assign w509[45] = |(datain[131:128] ^ 10);
  assign w509[46] = |(datain[127:124] ^ 0);
  assign w509[47] = |(datain[123:120] ^ 0);
  assign w509[48] = |(datain[119:116] ^ 0);
  assign w509[49] = |(datain[115:112] ^ 0);
  assign w509[50] = |(datain[111:108] ^ 12);
  assign w509[51] = |(datain[107:104] ^ 13);
  assign w509[52] = |(datain[103:100] ^ 2);
  assign w509[53] = |(datain[99:96] ^ 1);
  assign w509[54] = |(datain[95:92] ^ 11);
  assign w509[55] = |(datain[91:88] ^ 4);
  assign w509[56] = |(datain[87:84] ^ 4);
  assign w509[57] = |(datain[83:80] ^ 0);
  assign w509[58] = |(datain[79:76] ^ 8);
  assign w509[59] = |(datain[75:72] ^ 11);
  assign w509[60] = |(datain[71:68] ^ 9);
  assign w509[61] = |(datain[67:64] ^ 12);
  assign w509[62] = |(datain[63:60] ^ 6);
  assign w509[63] = |(datain[59:56] ^ 2);
  assign w509[64] = |(datain[55:52] ^ 0);
  assign w509[65] = |(datain[51:48] ^ 6);
  assign w509[66] = |(datain[47:44] ^ 11);
  assign w509[67] = |(datain[43:40] ^ 9);
  assign w509[68] = |(datain[39:36] ^ 2);
  assign w509[69] = |(datain[35:32] ^ 0);
  assign w509[70] = |(datain[31:28] ^ 0);
  assign w509[71] = |(datain[27:24] ^ 0);
  assign comp[509] = ~(|w509);
  wire [76-1:0] w510;
  assign w510[0] = |(datain[311:308] ^ 6);
  assign w510[1] = |(datain[307:304] ^ 6);
  assign w510[2] = |(datain[303:300] ^ 0);
  assign w510[3] = |(datain[299:296] ^ 6);
  assign w510[4] = |(datain[295:292] ^ 11);
  assign w510[5] = |(datain[291:288] ^ 10);
  assign w510[6] = |(datain[287:284] ^ 0);
  assign w510[7] = |(datain[283:280] ^ 6);
  assign w510[8] = |(datain[279:276] ^ 0);
  assign w510[9] = |(datain[275:272] ^ 6);
  assign w510[10] = |(datain[271:268] ^ 0);
  assign w510[11] = |(datain[267:264] ^ 3);
  assign w510[12] = |(datain[263:260] ^ 13);
  assign w510[13] = |(datain[259:256] ^ 6);
  assign w510[14] = |(datain[255:252] ^ 11);
  assign w510[15] = |(datain[251:248] ^ 4);
  assign w510[16] = |(datain[247:244] ^ 1);
  assign w510[17] = |(datain[243:240] ^ 10);
  assign w510[18] = |(datain[239:236] ^ 12);
  assign w510[19] = |(datain[235:232] ^ 13);
  assign w510[20] = |(datain[231:228] ^ 2);
  assign w510[21] = |(datain[227:224] ^ 1);
  assign w510[22] = |(datain[223:220] ^ 11);
  assign w510[23] = |(datain[219:216] ^ 10);
  assign w510[24] = |(datain[215:212] ^ 6);
  assign w510[25] = |(datain[211:208] ^ 10);
  assign w510[26] = |(datain[207:204] ^ 0);
  assign w510[27] = |(datain[203:200] ^ 6);
  assign w510[28] = |(datain[199:196] ^ 0);
  assign w510[29] = |(datain[195:192] ^ 3);
  assign w510[30] = |(datain[191:188] ^ 13);
  assign w510[31] = |(datain[187:184] ^ 6);
  assign w510[32] = |(datain[183:180] ^ 11);
  assign w510[33] = |(datain[179:176] ^ 4);
  assign w510[34] = |(datain[175:172] ^ 4);
  assign w510[35] = |(datain[171:168] ^ 14);
  assign w510[36] = |(datain[167:164] ^ 3);
  assign w510[37] = |(datain[163:160] ^ 3);
  assign w510[38] = |(datain[159:156] ^ 12);
  assign w510[39] = |(datain[155:152] ^ 9);
  assign w510[40] = |(datain[151:148] ^ 11);
  assign w510[41] = |(datain[147:144] ^ 1);
  assign w510[42] = |(datain[143:140] ^ 2);
  assign w510[43] = |(datain[139:136] ^ 7);
  assign w510[44] = |(datain[135:132] ^ 12);
  assign w510[45] = |(datain[131:128] ^ 13);
  assign w510[46] = |(datain[127:124] ^ 2);
  assign w510[47] = |(datain[123:120] ^ 1);
  assign w510[48] = |(datain[119:116] ^ 7);
  assign w510[49] = |(datain[115:112] ^ 2);
  assign w510[50] = |(datain[111:108] ^ 0);
  assign w510[51] = |(datain[107:104] ^ 7);
  assign w510[52] = |(datain[103:100] ^ 14);
  assign w510[53] = |(datain[99:96] ^ 8);
  assign w510[54] = |(datain[95:92] ^ 1);
  assign w510[55] = |(datain[91:88] ^ 3);
  assign w510[56] = |(datain[87:84] ^ 15);
  assign w510[57] = |(datain[83:80] ^ 15);
  assign w510[58] = |(datain[79:76] ^ 11);
  assign w510[59] = |(datain[75:72] ^ 4);
  assign w510[60] = |(datain[71:68] ^ 4);
  assign w510[61] = |(datain[67:64] ^ 15);
  assign w510[62] = |(datain[63:60] ^ 14);
  assign w510[63] = |(datain[59:56] ^ 11);
  assign w510[64] = |(datain[55:52] ^ 15);
  assign w510[65] = |(datain[51:48] ^ 1);
  assign w510[66] = |(datain[47:44] ^ 1);
  assign w510[67] = |(datain[43:40] ^ 14);
  assign w510[68] = |(datain[39:36] ^ 8);
  assign w510[69] = |(datain[35:32] ^ 11);
  assign w510[70] = |(datain[31:28] ^ 9);
  assign w510[71] = |(datain[27:24] ^ 4);
  assign w510[72] = |(datain[23:20] ^ 6);
  assign w510[73] = |(datain[19:16] ^ 8);
  assign w510[74] = |(datain[15:12] ^ 0);
  assign w510[75] = |(datain[11:8] ^ 6);
  assign comp[510] = ~(|w510);
  wire [50-1:0] w511;
  assign w511[0] = |(datain[311:308] ^ 2);
  assign w511[1] = |(datain[307:304] ^ 1);
  assign w511[2] = |(datain[303:300] ^ 12);
  assign w511[3] = |(datain[299:296] ^ 13);
  assign w511[4] = |(datain[295:292] ^ 12);
  assign w511[5] = |(datain[291:288] ^ 13);
  assign w511[6] = |(datain[287:284] ^ 8);
  assign w511[7] = |(datain[283:280] ^ 7);
  assign w511[8] = |(datain[279:276] ^ 13);
  assign w511[9] = |(datain[275:272] ^ 1);
  assign w511[10] = |(datain[271:268] ^ 11);
  assign w511[11] = |(datain[267:264] ^ 15);
  assign w511[12] = |(datain[263:260] ^ 0);
  assign w511[13] = |(datain[259:256] ^ 0);
  assign w511[14] = |(datain[255:252] ^ 0);
  assign w511[15] = |(datain[251:248] ^ 1);
  assign w511[16] = |(datain[247:244] ^ 15);
  assign w511[17] = |(datain[243:240] ^ 3);
  assign w511[18] = |(datain[239:236] ^ 10);
  assign w511[19] = |(datain[235:232] ^ 10);
  assign w511[20] = |(datain[231:228] ^ 5);
  assign w511[21] = |(datain[227:224] ^ 4);
  assign w511[22] = |(datain[223:220] ^ 4);
  assign w511[23] = |(datain[219:216] ^ 8);
  assign w511[24] = |(datain[215:212] ^ 4);
  assign w511[25] = |(datain[211:208] ^ 5);
  assign w511[26] = |(datain[207:204] ^ 2);
  assign w511[27] = |(datain[203:200] ^ 0);
  assign w511[28] = |(datain[199:196] ^ 4);
  assign w511[29] = |(datain[195:192] ^ 1);
  assign w511[30] = |(datain[191:188] ^ 5);
  assign w511[31] = |(datain[187:184] ^ 0);
  assign w511[32] = |(datain[183:180] ^ 5);
  assign w511[33] = |(datain[179:176] ^ 0);
  assign w511[34] = |(datain[175:172] ^ 4);
  assign w511[35] = |(datain[171:168] ^ 1);
  assign w511[36] = |(datain[167:164] ^ 5);
  assign w511[37] = |(datain[163:160] ^ 2);
  assign w511[38] = |(datain[159:156] ^ 4);
  assign w511[39] = |(datain[155:152] ^ 9);
  assign w511[40] = |(datain[151:148] ^ 5);
  assign w511[41] = |(datain[147:144] ^ 4);
  assign w511[42] = |(datain[143:140] ^ 4);
  assign w511[43] = |(datain[139:136] ^ 9);
  assign w511[44] = |(datain[135:132] ^ 4);
  assign w511[45] = |(datain[131:128] ^ 15);
  assign w511[46] = |(datain[127:124] ^ 4);
  assign w511[47] = |(datain[123:120] ^ 14);
  assign w511[48] = |(datain[119:116] ^ 0);
  assign w511[49] = |(datain[115:112] ^ 0);
  assign comp[511] = ~(|w511);
  wire [30-1:0] w512;
  assign w512[0] = |(datain[311:308] ^ 15);
  assign w512[1] = |(datain[307:304] ^ 12);
  assign w512[2] = |(datain[303:300] ^ 4);
  assign w512[3] = |(datain[299:296] ^ 13);
  assign w512[4] = |(datain[295:292] ^ 5);
  assign w512[5] = |(datain[291:288] ^ 10);
  assign w512[6] = |(datain[287:284] ^ 7);
  assign w512[7] = |(datain[283:280] ^ 5);
  assign w512[8] = |(datain[279:276] ^ 1);
  assign w512[9] = |(datain[275:272] ^ 13);
  assign w512[10] = |(datain[271:268] ^ 1);
  assign w512[11] = |(datain[267:264] ^ 15);
  assign w512[12] = |(datain[263:260] ^ 2);
  assign w512[13] = |(datain[259:256] ^ 14);
  assign w512[14] = |(datain[255:252] ^ 8);
  assign w512[15] = |(datain[251:248] ^ 11);
  assign w512[16] = |(datain[247:244] ^ 8);
  assign w512[17] = |(datain[243:240] ^ 4);
  assign w512[18] = |(datain[239:236] ^ 11);
  assign w512[19] = |(datain[235:232] ^ 11);
  assign w512[20] = |(datain[231:228] ^ 15);
  assign w512[21] = |(datain[227:224] ^ 12);
  assign w512[22] = |(datain[223:220] ^ 2);
  assign w512[23] = |(datain[219:216] ^ 14);
  assign w512[24] = |(datain[215:212] ^ 8);
  assign w512[25] = |(datain[211:208] ^ 11);
  assign w512[26] = |(datain[207:204] ^ 9);
  assign w512[27] = |(datain[203:200] ^ 12);
  assign w512[28] = |(datain[199:196] ^ 11);
  assign w512[29] = |(datain[195:192] ^ 9);
  assign comp[512] = ~(|w512);
  wire [30-1:0] w513;
  assign w513[0] = |(datain[311:308] ^ 8);
  assign w513[1] = |(datain[307:304] ^ 1);
  assign w513[2] = |(datain[303:300] ^ 0);
  assign w513[3] = |(datain[299:296] ^ 4);
  assign w513[4] = |(datain[295:292] ^ 11);
  assign w513[5] = |(datain[291:288] ^ 9);
  assign w513[6] = |(datain[287:284] ^ 0);
  assign w513[7] = |(datain[283:280] ^ 0);
  assign w513[8] = |(datain[279:276] ^ 15);
  assign w513[9] = |(datain[275:272] ^ 15);
  assign w513[10] = |(datain[271:268] ^ 8);
  assign w513[11] = |(datain[267:264] ^ 1);
  assign w513[12] = |(datain[263:260] ^ 14);
  assign w513[13] = |(datain[259:256] ^ 9);
  assign w513[14] = |(datain[255:252] ^ 8);
  assign w513[15] = |(datain[251:248] ^ 1);
  assign w513[16] = |(datain[247:244] ^ 0);
  assign w513[17] = |(datain[243:240] ^ 4);
  assign w513[18] = |(datain[239:236] ^ 11);
  assign w513[19] = |(datain[235:232] ^ 4);
  assign w513[20] = |(datain[231:228] ^ 13);
  assign w513[21] = |(datain[227:224] ^ 13);
  assign w513[22] = |(datain[223:220] ^ 12);
  assign w513[23] = |(datain[219:216] ^ 13);
  assign w513[24] = |(datain[215:212] ^ 2);
  assign w513[25] = |(datain[211:208] ^ 1);
  assign w513[26] = |(datain[207:204] ^ 14);
  assign w513[27] = |(datain[203:200] ^ 11);
  assign w513[28] = |(datain[199:196] ^ 2);
  assign w513[29] = |(datain[195:192] ^ 3);
  assign comp[513] = ~(|w513);
  wire [30-1:0] w514;
  assign w514[0] = |(datain[311:308] ^ 1);
  assign w514[1] = |(datain[307:304] ^ 14);
  assign w514[2] = |(datain[303:300] ^ 2);
  assign w514[3] = |(datain[299:296] ^ 5);
  assign w514[4] = |(datain[295:292] ^ 0);
  assign w514[5] = |(datain[291:288] ^ 0);
  assign w514[6] = |(datain[287:284] ^ 0);
  assign w514[7] = |(datain[283:280] ^ 11);
  assign w514[8] = |(datain[279:276] ^ 13);
  assign w514[9] = |(datain[275:272] ^ 11);
  assign w514[10] = |(datain[271:268] ^ 7);
  assign w514[11] = |(datain[267:264] ^ 4);
  assign w514[12] = |(datain[263:260] ^ 1);
  assign w514[13] = |(datain[259:256] ^ 3);
  assign w514[14] = |(datain[255:252] ^ 11);
  assign w514[15] = |(datain[251:248] ^ 9);
  assign w514[16] = |(datain[247:244] ^ 0);
  assign w514[17] = |(datain[243:240] ^ 0);
  assign w514[18] = |(datain[239:236] ^ 8);
  assign w514[19] = |(datain[235:232] ^ 0);
  assign w514[20] = |(datain[231:228] ^ 15);
  assign w514[21] = |(datain[227:224] ^ 3);
  assign w514[22] = |(datain[223:220] ^ 10);
  assign w514[23] = |(datain[219:216] ^ 5);
  assign w514[24] = |(datain[215:212] ^ 0);
  assign w514[25] = |(datain[211:208] ^ 5);
  assign w514[26] = |(datain[207:204] ^ 0);
  assign w514[27] = |(datain[203:200] ^ 0);
  assign w514[28] = |(datain[199:196] ^ 1);
  assign w514[29] = |(datain[195:192] ^ 0);
  assign comp[514] = ~(|w514);
  wire [28-1:0] w515;
  assign w515[0] = |(datain[311:308] ^ 8);
  assign w515[1] = |(datain[307:304] ^ 12);
  assign w515[2] = |(datain[303:300] ^ 0);
  assign w515[3] = |(datain[299:296] ^ 6);
  assign w515[4] = |(datain[295:292] ^ 2);
  assign w515[5] = |(datain[291:288] ^ 11);
  assign w515[6] = |(datain[287:284] ^ 0);
  assign w515[7] = |(datain[283:280] ^ 0);
  assign w515[8] = |(datain[279:276] ^ 11);
  assign w515[9] = |(datain[275:272] ^ 8);
  assign w515[10] = |(datain[271:268] ^ 2);
  assign w515[11] = |(datain[267:264] ^ 1);
  assign w515[12] = |(datain[263:260] ^ 3);
  assign w515[13] = |(datain[259:256] ^ 5);
  assign w515[14] = |(datain[255:252] ^ 12);
  assign w515[15] = |(datain[251:248] ^ 13);
  assign w515[16] = |(datain[247:244] ^ 2);
  assign w515[17] = |(datain[243:240] ^ 1);
  assign w515[18] = |(datain[239:236] ^ 8);
  assign w515[19] = |(datain[235:232] ^ 9);
  assign w515[20] = |(datain[231:228] ^ 1);
  assign w515[21] = |(datain[227:224] ^ 14);
  assign w515[22] = |(datain[223:220] ^ 0);
  assign w515[23] = |(datain[219:216] ^ 15);
  assign w515[24] = |(datain[215:212] ^ 0);
  assign w515[25] = |(datain[211:208] ^ 0);
  assign w515[26] = |(datain[207:204] ^ 8);
  assign w515[27] = |(datain[203:200] ^ 12);
  assign comp[515] = ~(|w515);
  wire [76-1:0] w516;
  assign w516[0] = |(datain[311:308] ^ 3);
  assign w516[1] = |(datain[307:304] ^ 4);
  assign w516[2] = |(datain[303:300] ^ 0);
  assign w516[3] = |(datain[299:296] ^ 1);
  assign w516[4] = |(datain[295:292] ^ 11);
  assign w516[5] = |(datain[291:288] ^ 4);
  assign w516[6] = |(datain[287:284] ^ 1);
  assign w516[7] = |(datain[283:280] ^ 9);
  assign w516[8] = |(datain[279:276] ^ 12);
  assign w516[9] = |(datain[275:272] ^ 13);
  assign w516[10] = |(datain[271:268] ^ 2);
  assign w516[11] = |(datain[267:264] ^ 1);
  assign w516[12] = |(datain[263:260] ^ 0);
  assign w516[13] = |(datain[259:256] ^ 4);
  assign w516[14] = |(datain[255:252] ^ 4);
  assign w516[15] = |(datain[251:248] ^ 1);
  assign w516[16] = |(datain[247:244] ^ 2);
  assign w516[17] = |(datain[243:240] ^ 14);
  assign w516[18] = |(datain[239:236] ^ 10);
  assign w516[19] = |(datain[235:232] ^ 2);
  assign w516[20] = |(datain[231:228] ^ 6);
  assign w516[21] = |(datain[227:224] ^ 5);
  assign w516[22] = |(datain[223:220] ^ 0);
  assign w516[23] = |(datain[219:216] ^ 3);
  assign w516[24] = |(datain[215:212] ^ 2);
  assign w516[25] = |(datain[211:208] ^ 14);
  assign w516[26] = |(datain[207:204] ^ 10);
  assign w516[27] = |(datain[203:200] ^ 2);
  assign w516[28] = |(datain[199:196] ^ 11);
  assign w516[29] = |(datain[195:192] ^ 1);
  assign w516[30] = |(datain[191:188] ^ 0);
  assign w516[31] = |(datain[187:184] ^ 3);
  assign w516[32] = |(datain[183:180] ^ 11);
  assign w516[33] = |(datain[179:176] ^ 15);
  assign w516[34] = |(datain[175:172] ^ 6);
  assign w516[35] = |(datain[171:168] ^ 7);
  assign w516[36] = |(datain[167:164] ^ 0);
  assign w516[37] = |(datain[163:160] ^ 3);
  assign w516[38] = |(datain[159:156] ^ 5);
  assign w516[39] = |(datain[155:152] ^ 7);
  assign w516[40] = |(datain[151:148] ^ 8);
  assign w516[41] = |(datain[147:144] ^ 11);
  assign w516[42] = |(datain[143:140] ^ 15);
  assign w516[43] = |(datain[139:136] ^ 2);
  assign w516[44] = |(datain[135:132] ^ 8);
  assign w516[45] = |(datain[131:128] ^ 0);
  assign w516[46] = |(datain[127:124] ^ 7);
  assign w516[47] = |(datain[123:120] ^ 12);
  assign w516[48] = |(datain[119:116] ^ 0);
  assign w516[49] = |(datain[115:112] ^ 1);
  assign w516[50] = |(datain[111:108] ^ 3);
  assign w516[51] = |(datain[107:104] ^ 10);
  assign w516[52] = |(datain[103:100] ^ 7);
  assign w516[53] = |(datain[99:96] ^ 5);
  assign w516[54] = |(datain[95:92] ^ 0);
  assign w516[55] = |(datain[91:88] ^ 13);
  assign w516[56] = |(datain[87:84] ^ 8);
  assign w516[57] = |(datain[83:80] ^ 10);
  assign w516[58] = |(datain[79:76] ^ 0);
  assign w516[59] = |(datain[75:72] ^ 4);
  assign w516[60] = |(datain[71:68] ^ 2);
  assign w516[61] = |(datain[67:64] ^ 14);
  assign w516[62] = |(datain[63:60] ^ 10);
  assign w516[63] = |(datain[59:56] ^ 2);
  assign w516[64] = |(datain[55:52] ^ 6);
  assign w516[65] = |(datain[51:48] ^ 5);
  assign w516[66] = |(datain[47:44] ^ 0);
  assign w516[67] = |(datain[43:40] ^ 3);
  assign w516[68] = |(datain[39:36] ^ 2);
  assign w516[69] = |(datain[35:32] ^ 14);
  assign w516[70] = |(datain[31:28] ^ 10);
  assign w516[71] = |(datain[27:24] ^ 2);
  assign w516[72] = |(datain[23:20] ^ 11);
  assign w516[73] = |(datain[19:16] ^ 1);
  assign w516[74] = |(datain[15:12] ^ 0);
  assign w516[75] = |(datain[11:8] ^ 3);
  assign comp[516] = ~(|w516);
  wire [60-1:0] w517;
  assign w517[0] = |(datain[311:308] ^ 1);
  assign w517[1] = |(datain[307:304] ^ 7);
  assign w517[2] = |(datain[303:300] ^ 0);
  assign w517[3] = |(datain[299:296] ^ 0);
  assign w517[4] = |(datain[295:292] ^ 11);
  assign w517[5] = |(datain[291:288] ^ 11);
  assign w517[6] = |(datain[287:284] ^ 1);
  assign w517[7] = |(datain[283:280] ^ 7);
  assign w517[8] = |(datain[279:276] ^ 0);
  assign w517[9] = |(datain[275:272] ^ 0);
  assign w517[10] = |(datain[271:268] ^ 0);
  assign w517[11] = |(datain[267:264] ^ 14);
  assign w517[12] = |(datain[263:260] ^ 1);
  assign w517[13] = |(datain[259:256] ^ 15);
  assign w517[14] = |(datain[255:252] ^ 11);
  assign w517[15] = |(datain[251:248] ^ 4);
  assign w517[16] = |(datain[247:244] ^ 13);
  assign w517[17] = |(datain[243:240] ^ 14);
  assign w517[18] = |(datain[239:236] ^ 12);
  assign w517[19] = |(datain[235:232] ^ 13);
  assign w517[20] = |(datain[231:228] ^ 2);
  assign w517[21] = |(datain[227:224] ^ 1);
  assign w517[22] = |(datain[223:220] ^ 11);
  assign w517[23] = |(datain[219:216] ^ 4);
  assign w517[24] = |(datain[215:212] ^ 2);
  assign w517[25] = |(datain[211:208] ^ 10);
  assign w517[26] = |(datain[207:204] ^ 12);
  assign w517[27] = |(datain[203:200] ^ 13);
  assign w517[28] = |(datain[199:196] ^ 2);
  assign w517[29] = |(datain[195:192] ^ 1);
  assign w517[30] = |(datain[191:188] ^ 8);
  assign w517[31] = |(datain[187:184] ^ 1);
  assign w517[32] = |(datain[183:180] ^ 15);
  assign w517[33] = |(datain[179:176] ^ 10);
  assign w517[34] = |(datain[175:172] ^ 0);
  assign w517[35] = |(datain[171:168] ^ 1);
  assign w517[36] = |(datain[167:164] ^ 0);
  assign w517[37] = |(datain[163:160] ^ 4);
  assign w517[38] = |(datain[159:156] ^ 7);
  assign w517[39] = |(datain[155:152] ^ 4);
  assign w517[40] = |(datain[151:148] ^ 2);
  assign w517[41] = |(datain[147:144] ^ 2);
  assign w517[42] = |(datain[143:140] ^ 8);
  assign w517[43] = |(datain[139:136] ^ 1);
  assign w517[44] = |(datain[135:132] ^ 15);
  assign w517[45] = |(datain[131:128] ^ 9);
  assign w517[46] = |(datain[127:124] ^ 11);
  assign w517[47] = |(datain[123:120] ^ 12);
  assign w517[48] = |(datain[119:116] ^ 0);
  assign w517[49] = |(datain[115:112] ^ 7);
  assign w517[50] = |(datain[111:108] ^ 7);
  assign w517[51] = |(datain[107:104] ^ 5);
  assign w517[52] = |(datain[103:100] ^ 0);
  assign w517[53] = |(datain[99:96] ^ 6);
  assign w517[54] = |(datain[95:92] ^ 14);
  assign w517[55] = |(datain[91:88] ^ 8);
  assign w517[56] = |(datain[87:84] ^ 12);
  assign w517[57] = |(datain[83:80] ^ 5);
  assign w517[58] = |(datain[79:76] ^ 0);
  assign w517[59] = |(datain[75:72] ^ 4);
  assign comp[517] = ~(|w517);
  wire [54-1:0] w518;
  assign w518[0] = |(datain[311:308] ^ 0);
  assign w518[1] = |(datain[307:304] ^ 1);
  assign w518[2] = |(datain[303:300] ^ 0);
  assign w518[3] = |(datain[299:296] ^ 0);
  assign w518[4] = |(datain[295:292] ^ 4);
  assign w518[5] = |(datain[291:288] ^ 14);
  assign w518[6] = |(datain[287:284] ^ 5);
  assign w518[7] = |(datain[283:280] ^ 0);
  assign w518[8] = |(datain[279:276] ^ 14);
  assign w518[9] = |(datain[275:272] ^ 8);
  assign w518[10] = |(datain[271:268] ^ 0);
  assign w518[11] = |(datain[267:264] ^ 0);
  assign w518[12] = |(datain[263:260] ^ 0);
  assign w518[13] = |(datain[259:256] ^ 0);
  assign w518[14] = |(datain[255:252] ^ 5);
  assign w518[15] = |(datain[251:248] ^ 13);
  assign w518[16] = |(datain[247:244] ^ 8);
  assign w518[17] = |(datain[243:240] ^ 1);
  assign w518[18] = |(datain[239:236] ^ 14);
  assign w518[19] = |(datain[235:232] ^ 13);
  assign w518[20] = |(datain[231:228] ^ 0);
  assign w518[21] = |(datain[227:224] ^ 8);
  assign w518[22] = |(datain[223:220] ^ 0);
  assign w518[23] = |(datain[219:216] ^ 1);
  assign w518[24] = |(datain[215:212] ^ 8);
  assign w518[25] = |(datain[211:208] ^ 13);
  assign w518[26] = |(datain[207:204] ^ 11);
  assign w518[27] = |(datain[203:200] ^ 6);
  assign w518[28] = |(datain[199:196] ^ 1);
  assign w518[29] = |(datain[195:192] ^ 12);
  assign w518[30] = |(datain[191:188] ^ 0);
  assign w518[31] = |(datain[187:184] ^ 1);
  assign w518[32] = |(datain[183:180] ^ 8);
  assign w518[33] = |(datain[179:176] ^ 9);
  assign w518[34] = |(datain[175:172] ^ 15);
  assign w518[35] = |(datain[171:168] ^ 7);
  assign w518[36] = |(datain[167:164] ^ 11);
  assign w518[37] = |(datain[163:160] ^ 9);
  assign w518[38] = |(datain[159:156] ^ 8);
  assign w518[39] = |(datain[155:152] ^ 11);
  assign w518[40] = |(datain[151:148] ^ 0);
  assign w518[41] = |(datain[147:144] ^ 1);
  assign w518[42] = |(datain[143:140] ^ 10);
  assign w518[43] = |(datain[139:136] ^ 12);
  assign w518[44] = |(datain[135:132] ^ 0);
  assign w518[45] = |(datain[131:128] ^ 4);
  assign w518[46] = |(datain[127:124] ^ 0);
  assign w518[47] = |(datain[123:120] ^ 0);
  assign w518[48] = |(datain[119:116] ^ 10);
  assign w518[49] = |(datain[115:112] ^ 10);
  assign w518[50] = |(datain[111:108] ^ 14);
  assign w518[51] = |(datain[107:104] ^ 2);
  assign w518[52] = |(datain[103:100] ^ 15);
  assign w518[53] = |(datain[99:96] ^ 10);
  assign comp[518] = ~(|w518);
  wire [46-1:0] w519;
  assign w519[0] = |(datain[311:308] ^ 14);
  assign w519[1] = |(datain[307:304] ^ 8);
  assign w519[2] = |(datain[303:300] ^ 0);
  assign w519[3] = |(datain[299:296] ^ 0);
  assign w519[4] = |(datain[295:292] ^ 0);
  assign w519[5] = |(datain[291:288] ^ 0);
  assign w519[6] = |(datain[287:284] ^ 5);
  assign w519[7] = |(datain[283:280] ^ 13);
  assign w519[8] = |(datain[279:276] ^ 8);
  assign w519[9] = |(datain[275:272] ^ 1);
  assign w519[10] = |(datain[271:268] ^ 14);
  assign w519[11] = |(datain[267:264] ^ 13);
  assign w519[12] = |(datain[263:260] ^ 0);
  assign w519[13] = |(datain[259:256] ^ 8);
  assign w519[14] = |(datain[255:252] ^ 0);
  assign w519[15] = |(datain[251:248] ^ 1);
  assign w519[16] = |(datain[247:244] ^ 8);
  assign w519[17] = |(datain[243:240] ^ 13);
  assign w519[18] = |(datain[239:236] ^ 11);
  assign w519[19] = |(datain[235:232] ^ 6);
  assign w519[20] = |(datain[231:228] ^ 1);
  assign w519[21] = |(datain[227:224] ^ 12);
  assign w519[22] = |(datain[223:220] ^ 0);
  assign w519[23] = |(datain[219:216] ^ 1);
  assign w519[24] = |(datain[215:212] ^ 8);
  assign w519[25] = |(datain[211:208] ^ 11);
  assign w519[26] = |(datain[207:204] ^ 15);
  assign w519[27] = |(datain[203:200] ^ 14);
  assign w519[28] = |(datain[199:196] ^ 11);
  assign w519[29] = |(datain[195:192] ^ 9);
  assign w519[30] = |(datain[191:188] ^ 8);
  assign w519[31] = |(datain[187:184] ^ 11);
  assign w519[32] = |(datain[183:180] ^ 0);
  assign w519[33] = |(datain[179:176] ^ 1);
  assign w519[34] = |(datain[175:172] ^ 10);
  assign w519[35] = |(datain[171:168] ^ 12);
  assign w519[36] = |(datain[167:164] ^ 0);
  assign w519[37] = |(datain[163:160] ^ 4);
  assign w519[38] = |(datain[159:156] ^ 0);
  assign w519[39] = |(datain[155:152] ^ 0);
  assign w519[40] = |(datain[151:148] ^ 10);
  assign w519[41] = |(datain[147:144] ^ 10);
  assign w519[42] = |(datain[143:140] ^ 14);
  assign w519[43] = |(datain[139:136] ^ 2);
  assign w519[44] = |(datain[135:132] ^ 15);
  assign w519[45] = |(datain[131:128] ^ 10);
  assign comp[519] = ~(|w519);
  wire [76-1:0] w520;
  assign w520[0] = |(datain[311:308] ^ 14);
  assign w520[1] = |(datain[307:304] ^ 9);
  assign w520[2] = |(datain[303:300] ^ 1);
  assign w520[3] = |(datain[299:296] ^ 15);
  assign w520[4] = |(datain[295:292] ^ 15);
  assign w520[5] = |(datain[291:288] ^ 15);
  assign w520[6] = |(datain[287:284] ^ 11);
  assign w520[7] = |(datain[283:280] ^ 8);
  assign w520[8] = |(datain[279:276] ^ 1);
  assign w520[9] = |(datain[275:272] ^ 0);
  assign w520[10] = |(datain[271:268] ^ 0);
  assign w520[11] = |(datain[267:264] ^ 5);
  assign w520[12] = |(datain[263:260] ^ 11);
  assign w520[13] = |(datain[259:256] ^ 10);
  assign w520[14] = |(datain[255:252] ^ 8);
  assign w520[15] = |(datain[251:248] ^ 0);
  assign w520[16] = |(datain[247:244] ^ 0);
  assign w520[17] = |(datain[243:240] ^ 0);
  assign w520[18] = |(datain[239:236] ^ 11);
  assign w520[19] = |(datain[235:232] ^ 9);
  assign w520[20] = |(datain[231:228] ^ 1);
  assign w520[21] = |(datain[227:224] ^ 0);
  assign w520[22] = |(datain[223:220] ^ 0);
  assign w520[23] = |(datain[219:216] ^ 0);
  assign w520[24] = |(datain[215:212] ^ 12);
  assign w520[25] = |(datain[211:208] ^ 13);
  assign w520[26] = |(datain[207:204] ^ 1);
  assign w520[27] = |(datain[203:200] ^ 3);
  assign w520[28] = |(datain[199:196] ^ 12);
  assign w520[29] = |(datain[195:192] ^ 15);
  assign w520[30] = |(datain[191:188] ^ 3);
  assign w520[31] = |(datain[187:184] ^ 2);
  assign w520[32] = |(datain[183:180] ^ 12);
  assign w520[33] = |(datain[179:176] ^ 0);
  assign w520[34] = |(datain[175:172] ^ 12);
  assign w520[35] = |(datain[171:168] ^ 15);
  assign w520[36] = |(datain[167:164] ^ 11);
  assign w520[37] = |(datain[163:160] ^ 4);
  assign w520[38] = |(datain[159:156] ^ 4);
  assign w520[39] = |(datain[155:152] ^ 0);
  assign w520[40] = |(datain[151:148] ^ 8);
  assign w520[41] = |(datain[147:144] ^ 13);
  assign w520[42] = |(datain[143:140] ^ 9);
  assign w520[43] = |(datain[139:136] ^ 6);
  assign w520[44] = |(datain[135:132] ^ 0);
  assign w520[45] = |(datain[131:128] ^ 0);
  assign w520[46] = |(datain[127:124] ^ 0);
  assign w520[47] = |(datain[123:120] ^ 1);
  assign w520[48] = |(datain[119:116] ^ 2);
  assign w520[49] = |(datain[115:112] ^ 14);
  assign w520[50] = |(datain[111:108] ^ 8);
  assign w520[51] = |(datain[107:104] ^ 11);
  assign w520[52] = |(datain[103:100] ^ 8);
  assign w520[53] = |(datain[99:96] ^ 14);
  assign w520[54] = |(datain[95:92] ^ 14);
  assign w520[55] = |(datain[91:88] ^ 13);
  assign w520[56] = |(datain[87:84] ^ 0);
  assign w520[57] = |(datain[83:80] ^ 3);
  assign w520[58] = |(datain[79:76] ^ 2);
  assign w520[59] = |(datain[75:72] ^ 14);
  assign w520[60] = |(datain[71:68] ^ 8);
  assign w520[61] = |(datain[67:64] ^ 11);
  assign w520[62] = |(datain[63:60] ^ 9);
  assign w520[63] = |(datain[59:56] ^ 14);
  assign w520[64] = |(datain[55:52] ^ 1);
  assign w520[65] = |(datain[51:48] ^ 11);
  assign w520[66] = |(datain[47:44] ^ 0);
  assign w520[67] = |(datain[43:40] ^ 1);
  assign w520[68] = |(datain[39:36] ^ 12);
  assign w520[69] = |(datain[35:32] ^ 13);
  assign w520[70] = |(datain[31:28] ^ 2);
  assign w520[71] = |(datain[27:24] ^ 1);
  assign w520[72] = |(datain[23:20] ^ 3);
  assign w520[73] = |(datain[19:16] ^ 11);
  assign w520[74] = |(datain[15:12] ^ 12);
  assign w520[75] = |(datain[11:8] ^ 1);
  assign comp[520] = ~(|w520);
  wire [46-1:0] w521;
  assign w521[0] = |(datain[311:308] ^ 0);
  assign w521[1] = |(datain[307:304] ^ 14);
  assign w521[2] = |(datain[303:300] ^ 1);
  assign w521[3] = |(datain[299:296] ^ 15);
  assign w521[4] = |(datain[295:292] ^ 11);
  assign w521[5] = |(datain[291:288] ^ 14);
  assign w521[6] = |(datain[287:284] ^ 0);
  assign w521[7] = |(datain[283:280] ^ 3);
  assign w521[8] = |(datain[279:276] ^ 0);
  assign w521[9] = |(datain[275:272] ^ 1);
  assign w521[10] = |(datain[271:268] ^ 11);
  assign w521[11] = |(datain[267:264] ^ 10);
  assign w521[12] = |(datain[263:260] ^ 9);
  assign w521[13] = |(datain[259:256] ^ 6);
  assign w521[14] = |(datain[255:252] ^ 2);
  assign w521[15] = |(datain[251:248] ^ 7);
  assign w521[16] = |(datain[247:244] ^ 11);
  assign w521[17] = |(datain[243:240] ^ 9);
  assign w521[18] = |(datain[239:236] ^ 12);
  assign w521[19] = |(datain[235:232] ^ 1);
  assign w521[20] = |(datain[231:228] ^ 0);
  assign w521[21] = |(datain[227:224] ^ 2);
  assign w521[22] = |(datain[223:220] ^ 10);
  assign w521[23] = |(datain[219:216] ^ 12);
  assign w521[24] = |(datain[215:212] ^ 3);
  assign w521[25] = |(datain[211:208] ^ 2);
  assign w521[26] = |(datain[207:204] ^ 12);
  assign w521[27] = |(datain[203:200] ^ 2);
  assign w521[28] = |(datain[199:196] ^ 3);
  assign w521[29] = |(datain[195:192] ^ 2);
  assign w521[30] = |(datain[191:188] ^ 12);
  assign w521[31] = |(datain[187:184] ^ 6);
  assign w521[32] = |(datain[183:180] ^ 3);
  assign w521[33] = |(datain[179:176] ^ 2);
  assign w521[34] = |(datain[175:172] ^ 12);
  assign w521[35] = |(datain[171:168] ^ 1);
  assign w521[36] = |(datain[167:164] ^ 8);
  assign w521[37] = |(datain[163:160] ^ 8);
  assign w521[38] = |(datain[159:156] ^ 4);
  assign w521[39] = |(datain[155:152] ^ 4);
  assign w521[40] = |(datain[151:148] ^ 15);
  assign w521[41] = |(datain[147:144] ^ 15);
  assign w521[42] = |(datain[143:140] ^ 14);
  assign w521[43] = |(datain[139:136] ^ 2);
  assign w521[44] = |(datain[135:132] ^ 15);
  assign w521[45] = |(datain[131:128] ^ 4);
  assign comp[521] = ~(|w521);
  wire [34-1:0] w522;
  assign w522[0] = |(datain[311:308] ^ 9);
  assign w522[1] = |(datain[307:304] ^ 6);
  assign w522[2] = |(datain[303:300] ^ 3);
  assign w522[3] = |(datain[299:296] ^ 5);
  assign w522[4] = |(datain[295:292] ^ 0);
  assign w522[5] = |(datain[291:288] ^ 2);
  assign w522[6] = |(datain[287:284] ^ 8);
  assign w522[7] = |(datain[283:280] ^ 13);
  assign w522[8] = |(datain[279:276] ^ 11);
  assign w522[9] = |(datain[275:272] ^ 6);
  assign w522[10] = |(datain[271:268] ^ 0);
  assign w522[11] = |(datain[267:264] ^ 15);
  assign w522[12] = |(datain[263:260] ^ 0);
  assign w522[13] = |(datain[259:256] ^ 0);
  assign w522[14] = |(datain[255:252] ^ 11);
  assign w522[15] = |(datain[251:248] ^ 9);
  assign w522[16] = |(datain[247:244] ^ 1);
  assign w522[17] = |(datain[243:240] ^ 0);
  assign w522[18] = |(datain[239:236] ^ 0);
  assign w522[19] = |(datain[235:232] ^ 1);
  assign w522[20] = |(datain[231:228] ^ 3);
  assign w522[21] = |(datain[227:224] ^ 1);
  assign w522[22] = |(datain[223:220] ^ 1);
  assign w522[23] = |(datain[219:216] ^ 4);
  assign w522[24] = |(datain[215:212] ^ 4);
  assign w522[25] = |(datain[211:208] ^ 6);
  assign w522[26] = |(datain[207:204] ^ 4);
  assign w522[27] = |(datain[203:200] ^ 6);
  assign w522[28] = |(datain[199:196] ^ 14);
  assign w522[29] = |(datain[195:192] ^ 2);
  assign w522[30] = |(datain[191:188] ^ 15);
  assign w522[31] = |(datain[187:184] ^ 10);
  assign w522[32] = |(datain[183:180] ^ 12);
  assign w522[33] = |(datain[179:176] ^ 3);
  assign comp[522] = ~(|w522);
  wire [34-1:0] w523;
  assign w523[0] = |(datain[311:308] ^ 9);
  assign w523[1] = |(datain[307:304] ^ 6);
  assign w523[2] = |(datain[303:300] ^ 11);
  assign w523[3] = |(datain[299:296] ^ 10);
  assign w523[4] = |(datain[295:292] ^ 0);
  assign w523[5] = |(datain[291:288] ^ 2);
  assign w523[6] = |(datain[287:284] ^ 8);
  assign w523[7] = |(datain[283:280] ^ 13);
  assign w523[8] = |(datain[279:276] ^ 11);
  assign w523[9] = |(datain[275:272] ^ 6);
  assign w523[10] = |(datain[271:268] ^ 1);
  assign w523[11] = |(datain[267:264] ^ 1);
  assign w523[12] = |(datain[263:260] ^ 0);
  assign w523[13] = |(datain[259:256] ^ 0);
  assign w523[14] = |(datain[255:252] ^ 11);
  assign w523[15] = |(datain[251:248] ^ 9);
  assign w523[16] = |(datain[247:244] ^ 5);
  assign w523[17] = |(datain[243:240] ^ 2);
  assign w523[18] = |(datain[239:236] ^ 0);
  assign w523[19] = |(datain[235:232] ^ 1);
  assign w523[20] = |(datain[231:228] ^ 3);
  assign w523[21] = |(datain[227:224] ^ 1);
  assign w523[22] = |(datain[223:220] ^ 1);
  assign w523[23] = |(datain[219:216] ^ 4);
  assign w523[24] = |(datain[215:212] ^ 4);
  assign w523[25] = |(datain[211:208] ^ 6);
  assign w523[26] = |(datain[207:204] ^ 4);
  assign w523[27] = |(datain[203:200] ^ 6);
  assign w523[28] = |(datain[199:196] ^ 14);
  assign w523[29] = |(datain[195:192] ^ 2);
  assign w523[30] = |(datain[191:188] ^ 15);
  assign w523[31] = |(datain[187:184] ^ 10);
  assign w523[32] = |(datain[183:180] ^ 12);
  assign w523[33] = |(datain[179:176] ^ 3);
  assign comp[523] = ~(|w523);
  wire [32-1:0] w524;
  assign w524[0] = |(datain[311:308] ^ 3);
  assign w524[1] = |(datain[307:304] ^ 13);
  assign w524[2] = |(datain[303:300] ^ 0);
  assign w524[3] = |(datain[299:296] ^ 0);
  assign w524[4] = |(datain[295:292] ^ 4);
  assign w524[5] = |(datain[291:288] ^ 11);
  assign w524[6] = |(datain[287:284] ^ 7);
  assign w524[7] = |(datain[283:280] ^ 5);
  assign w524[8] = |(datain[279:276] ^ 3);
  assign w524[9] = |(datain[275:272] ^ 6);
  assign w524[10] = |(datain[271:268] ^ 8);
  assign w524[11] = |(datain[267:264] ^ 11);
  assign w524[12] = |(datain[263:260] ^ 14);
  assign w524[13] = |(datain[259:256] ^ 12);
  assign w524[14] = |(datain[255:252] ^ 8);
  assign w524[15] = |(datain[251:248] ^ 11);
  assign w524[16] = |(datain[247:244] ^ 7);
  assign w524[17] = |(datain[243:240] ^ 6);
  assign w524[18] = |(datain[239:236] ^ 0);
  assign w524[19] = |(datain[235:232] ^ 0);
  assign w524[20] = |(datain[231:228] ^ 8);
  assign w524[21] = |(datain[227:224] ^ 11);
  assign w524[22] = |(datain[223:220] ^ 7);
  assign w524[23] = |(datain[219:216] ^ 14);
  assign w524[24] = |(datain[215:212] ^ 0);
  assign w524[25] = |(datain[211:208] ^ 2);
  assign w524[26] = |(datain[207:204] ^ 8);
  assign w524[27] = |(datain[203:200] ^ 12);
  assign w524[28] = |(datain[199:196] ^ 12);
  assign w524[29] = |(datain[195:192] ^ 9);
  assign w524[30] = |(datain[191:188] ^ 8);
  assign w524[31] = |(datain[187:184] ^ 14);
  assign comp[524] = ~(|w524);
  wire [44-1:0] w525;
  assign w525[0] = |(datain[311:308] ^ 0);
  assign w525[1] = |(datain[307:304] ^ 1);
  assign w525[2] = |(datain[303:300] ^ 3);
  assign w525[3] = |(datain[299:296] ^ 3);
  assign w525[4] = |(datain[295:292] ^ 12);
  assign w525[5] = |(datain[291:288] ^ 0);
  assign w525[6] = |(datain[287:284] ^ 8);
  assign w525[7] = |(datain[283:280] ^ 10);
  assign w525[8] = |(datain[279:276] ^ 2);
  assign w525[9] = |(datain[275:272] ^ 6);
  assign w525[10] = |(datain[271:268] ^ 5);
  assign w525[11] = |(datain[267:264] ^ 15);
  assign w525[12] = |(datain[263:260] ^ 0);
  assign w525[13] = |(datain[259:256] ^ 1);
  assign w525[14] = |(datain[255:252] ^ 8);
  assign w525[15] = |(datain[251:248] ^ 8);
  assign w525[16] = |(datain[247:244] ^ 2);
  assign w525[17] = |(datain[243:240] ^ 6);
  assign w525[18] = |(datain[239:236] ^ 1);
  assign w525[19] = |(datain[235:232] ^ 6);
  assign w525[20] = |(datain[231:228] ^ 0);
  assign w525[21] = |(datain[227:224] ^ 2);
  assign w525[22] = |(datain[223:220] ^ 3);
  assign w525[23] = |(datain[219:216] ^ 3);
  assign w525[24] = |(datain[215:212] ^ 12);
  assign w525[25] = |(datain[211:208] ^ 0);
  assign w525[26] = |(datain[207:204] ^ 8);
  assign w525[27] = |(datain[203:200] ^ 0);
  assign w525[28] = |(datain[199:196] ^ 3);
  assign w525[29] = |(datain[195:192] ^ 14);
  assign w525[30] = |(datain[191:188] ^ 1);
  assign w525[31] = |(datain[187:184] ^ 3);
  assign w525[32] = |(datain[183:180] ^ 0);
  assign w525[33] = |(datain[179:176] ^ 2);
  assign w525[34] = |(datain[175:172] ^ 0);
  assign w525[35] = |(datain[171:168] ^ 1);
  assign w525[36] = |(datain[167:164] ^ 7);
  assign w525[37] = |(datain[163:160] ^ 4);
  assign w525[38] = |(datain[159:156] ^ 2);
  assign w525[39] = |(datain[155:152] ^ 12);
  assign w525[40] = |(datain[151:148] ^ 11);
  assign w525[41] = |(datain[147:144] ^ 4);
  assign w525[42] = |(datain[143:140] ^ 3);
  assign w525[43] = |(datain[139:136] ^ 13);
  assign comp[525] = ~(|w525);
  wire [76-1:0] w526;
  assign w526[0] = |(datain[311:308] ^ 0);
  assign w526[1] = |(datain[307:304] ^ 3);
  assign w526[2] = |(datain[303:300] ^ 14);
  assign w526[3] = |(datain[299:296] ^ 9);
  assign w526[4] = |(datain[295:292] ^ 12);
  assign w526[5] = |(datain[291:288] ^ 0);
  assign w526[6] = |(datain[287:284] ^ 0);
  assign w526[7] = |(datain[283:280] ^ 0);
  assign w526[8] = |(datain[279:276] ^ 11);
  assign w526[9] = |(datain[275:272] ^ 8);
  assign w526[10] = |(datain[271:268] ^ 0);
  assign w526[11] = |(datain[267:264] ^ 0);
  assign w526[12] = |(datain[263:260] ^ 4);
  assign w526[13] = |(datain[259:256] ^ 3);
  assign w526[14] = |(datain[255:252] ^ 11);
  assign w526[15] = |(datain[251:248] ^ 10);
  assign w526[16] = |(datain[247:244] ^ 1);
  assign w526[17] = |(datain[243:240] ^ 14);
  assign w526[18] = |(datain[239:236] ^ 15);
  assign w526[19] = |(datain[235:232] ^ 13);
  assign w526[20] = |(datain[231:228] ^ 12);
  assign w526[21] = |(datain[227:224] ^ 13);
  assign w526[22] = |(datain[223:220] ^ 2);
  assign w526[23] = |(datain[219:216] ^ 1);
  assign w526[24] = |(datain[215:212] ^ 5);
  assign w526[25] = |(datain[211:208] ^ 1);
  assign w526[26] = |(datain[207:204] ^ 11);
  assign w526[27] = |(datain[203:200] ^ 8);
  assign w526[28] = |(datain[199:196] ^ 0);
  assign w526[29] = |(datain[195:192] ^ 1);
  assign w526[30] = |(datain[191:188] ^ 4);
  assign w526[31] = |(datain[187:184] ^ 3);
  assign w526[32] = |(datain[183:180] ^ 3);
  assign w526[33] = |(datain[179:176] ^ 3);
  assign w526[34] = |(datain[175:172] ^ 12);
  assign w526[35] = |(datain[171:168] ^ 9);
  assign w526[36] = |(datain[167:164] ^ 12);
  assign w526[37] = |(datain[163:160] ^ 13);
  assign w526[38] = |(datain[159:156] ^ 2);
  assign w526[39] = |(datain[155:152] ^ 1);
  assign w526[40] = |(datain[151:148] ^ 12);
  assign w526[41] = |(datain[147:144] ^ 12);
  assign w526[42] = |(datain[143:140] ^ 11);
  assign w526[43] = |(datain[139:136] ^ 8);
  assign w526[44] = |(datain[135:132] ^ 0);
  assign w526[45] = |(datain[131:128] ^ 2);
  assign w526[46] = |(datain[127:124] ^ 3);
  assign w526[47] = |(datain[123:120] ^ 13);
  assign w526[48] = |(datain[119:116] ^ 11);
  assign w526[49] = |(datain[115:112] ^ 10);
  assign w526[50] = |(datain[111:108] ^ 1);
  assign w526[51] = |(datain[107:104] ^ 14);
  assign w526[52] = |(datain[103:100] ^ 15);
  assign w526[53] = |(datain[99:96] ^ 13);
  assign w526[54] = |(datain[95:92] ^ 12);
  assign w526[55] = |(datain[91:88] ^ 13);
  assign w526[56] = |(datain[87:84] ^ 2);
  assign w526[57] = |(datain[83:80] ^ 1);
  assign w526[58] = |(datain[79:76] ^ 9);
  assign w526[59] = |(datain[75:72] ^ 3);
  assign w526[60] = |(datain[71:68] ^ 11);
  assign w526[61] = |(datain[67:64] ^ 8);
  assign w526[62] = |(datain[63:60] ^ 0);
  assign w526[63] = |(datain[59:56] ^ 0);
  assign w526[64] = |(datain[55:52] ^ 5);
  assign w526[65] = |(datain[51:48] ^ 7);
  assign w526[66] = |(datain[47:44] ^ 12);
  assign w526[67] = |(datain[43:40] ^ 13);
  assign w526[68] = |(datain[39:36] ^ 2);
  assign w526[69] = |(datain[35:32] ^ 1);
  assign w526[70] = |(datain[31:28] ^ 5);
  assign w526[71] = |(datain[27:24] ^ 1);
  assign w526[72] = |(datain[23:20] ^ 5);
  assign w526[73] = |(datain[19:16] ^ 2);
  assign w526[74] = |(datain[15:12] ^ 11);
  assign w526[75] = |(datain[11:8] ^ 4);
  assign comp[526] = ~(|w526);
  wire [72-1:0] w527;
  assign w527[0] = |(datain[311:308] ^ 8);
  assign w527[1] = |(datain[307:304] ^ 11);
  assign w527[2] = |(datain[303:300] ^ 0);
  assign w527[3] = |(datain[299:296] ^ 15);
  assign w527[4] = |(datain[295:292] ^ 8);
  assign w527[5] = |(datain[291:288] ^ 3);
  assign w527[6] = |(datain[287:284] ^ 14);
  assign w527[7] = |(datain[283:280] ^ 9);
  assign w527[8] = |(datain[279:276] ^ 0);
  assign w527[9] = |(datain[275:272] ^ 3);
  assign w527[10] = |(datain[271:268] ^ 8);
  assign w527[11] = |(datain[267:264] ^ 1);
  assign w527[12] = |(datain[263:260] ^ 12);
  assign w527[13] = |(datain[259:256] ^ 1);
  assign w527[14] = |(datain[255:252] ^ 10);
  assign w527[15] = |(datain[251:248] ^ 10);
  assign w527[16] = |(datain[247:244] ^ 0);
  assign w527[17] = |(datain[243:240] ^ 0);
  assign w527[18] = |(datain[239:236] ^ 8);
  assign w527[19] = |(datain[235:232] ^ 11);
  assign w527[20] = |(datain[231:228] ^ 13);
  assign w527[21] = |(datain[227:224] ^ 8);
  assign w527[22] = |(datain[223:220] ^ 8);
  assign w527[23] = |(datain[219:216] ^ 9);
  assign w527[24] = |(datain[215:212] ^ 4);
  assign w527[25] = |(datain[211:208] ^ 15);
  assign w527[26] = |(datain[207:204] ^ 0);
  assign w527[27] = |(datain[203:200] ^ 1);
  assign w527[28] = |(datain[199:196] ^ 5);
  assign w527[29] = |(datain[195:192] ^ 11);
  assign w527[30] = |(datain[191:188] ^ 5);
  assign w527[31] = |(datain[187:184] ^ 3);
  assign w527[32] = |(datain[183:180] ^ 8);
  assign w527[33] = |(datain[179:176] ^ 1);
  assign w527[34] = |(datain[175:172] ^ 14);
  assign w527[35] = |(datain[171:168] ^ 11);
  assign w527[36] = |(datain[167:164] ^ 10);
  assign w527[37] = |(datain[163:160] ^ 9);
  assign w527[38] = |(datain[159:156] ^ 0);
  assign w527[39] = |(datain[155:152] ^ 0);
  assign w527[40] = |(datain[151:148] ^ 8);
  assign w527[41] = |(datain[147:144] ^ 11);
  assign w527[42] = |(datain[143:140] ^ 1);
  assign w527[43] = |(datain[139:136] ^ 15);
  assign w527[44] = |(datain[135:132] ^ 11);
  assign w527[45] = |(datain[131:128] ^ 9);
  assign w527[46] = |(datain[127:124] ^ 0);
  assign w527[47] = |(datain[123:120] ^ 3);
  assign w527[48] = |(datain[119:116] ^ 0);
  assign w527[49] = |(datain[115:112] ^ 0);
  assign w527[50] = |(datain[111:108] ^ 11);
  assign w527[51] = |(datain[107:104] ^ 4);
  assign w527[52] = |(datain[103:100] ^ 4);
  assign w527[53] = |(datain[99:96] ^ 0);
  assign w527[54] = |(datain[95:92] ^ 5);
  assign w527[55] = |(datain[91:88] ^ 10);
  assign w527[56] = |(datain[87:84] ^ 5);
  assign w527[57] = |(datain[83:80] ^ 2);
  assign w527[58] = |(datain[79:76] ^ 8);
  assign w527[59] = |(datain[75:72] ^ 1);
  assign w527[60] = |(datain[71:68] ^ 14);
  assign w527[61] = |(datain[67:64] ^ 10);
  assign w527[62] = |(datain[63:60] ^ 11);
  assign w527[63] = |(datain[59:56] ^ 2);
  assign w527[64] = |(datain[55:52] ^ 0);
  assign w527[65] = |(datain[51:48] ^ 0);
  assign w527[66] = |(datain[47:44] ^ 12);
  assign w527[67] = |(datain[43:40] ^ 13);
  assign w527[68] = |(datain[39:36] ^ 2);
  assign w527[69] = |(datain[35:32] ^ 1);
  assign w527[70] = |(datain[31:28] ^ 5);
  assign w527[71] = |(datain[27:24] ^ 11);
  assign comp[527] = ~(|w527);
  wire [56-1:0] w528;
  assign w528[0] = |(datain[311:308] ^ 5);
  assign w528[1] = |(datain[307:304] ^ 15);
  assign w528[2] = |(datain[303:300] ^ 8);
  assign w528[3] = |(datain[299:296] ^ 1);
  assign w528[4] = |(datain[295:292] ^ 14);
  assign w528[5] = |(datain[291:288] ^ 15);
  assign w528[6] = |(datain[287:284] ^ 0);
  assign w528[7] = |(datain[283:280] ^ 7);
  assign w528[8] = |(datain[279:276] ^ 0);
  assign w528[9] = |(datain[275:272] ^ 1);
  assign w528[10] = |(datain[271:268] ^ 14);
  assign w528[11] = |(datain[267:264] ^ 8);
  assign w528[12] = |(datain[263:260] ^ 0);
  assign w528[13] = |(datain[259:256] ^ 2);
  assign w528[14] = |(datain[255:252] ^ 0);
  assign w528[15] = |(datain[251:248] ^ 0);
  assign w528[16] = |(datain[247:244] ^ 14);
  assign w528[17] = |(datain[243:240] ^ 11);
  assign w528[18] = |(datain[239:236] ^ 1);
  assign w528[19] = |(datain[235:232] ^ 2);
  assign w528[20] = |(datain[231:228] ^ 8);
  assign w528[21] = |(datain[227:224] ^ 13);
  assign w528[22] = |(datain[223:220] ^ 11);
  assign w528[23] = |(datain[219:216] ^ 5);
  assign w528[24] = |(datain[215:212] ^ 2);
  assign w528[25] = |(datain[211:208] ^ 3);
  assign w528[26] = |(datain[207:204] ^ 0);
  assign w528[27] = |(datain[203:200] ^ 1);
  assign w528[28] = |(datain[199:196] ^ 11);
  assign w528[29] = |(datain[195:192] ^ 9);
  assign w528[30] = |(datain[191:188] ^ 11);
  assign w528[31] = |(datain[187:184] ^ 6);
  assign w528[32] = |(datain[183:180] ^ 0);
  assign w528[33] = |(datain[179:176] ^ 3);
  assign w528[34] = |(datain[175:172] ^ 8);
  assign w528[35] = |(datain[171:168] ^ 12);
  assign w528[36] = |(datain[167:164] ^ 12);
  assign w528[37] = |(datain[163:160] ^ 8);
  assign w528[38] = |(datain[159:156] ^ 8);
  assign w528[39] = |(datain[155:152] ^ 14);
  assign w528[40] = |(datain[151:148] ^ 13);
  assign w528[41] = |(datain[147:144] ^ 8);
  assign w528[42] = |(datain[143:140] ^ 8);
  assign w528[43] = |(datain[139:136] ^ 0);
  assign w528[44] = |(datain[135:132] ^ 0);
  assign w528[45] = |(datain[131:128] ^ 4);
  assign w528[46] = |(datain[127:124] ^ 0);
  assign w528[47] = |(datain[123:120] ^ 1);
  assign w528[48] = |(datain[119:116] ^ 4);
  assign w528[49] = |(datain[115:112] ^ 6);
  assign w528[50] = |(datain[111:108] ^ 14);
  assign w528[51] = |(datain[107:104] ^ 2);
  assign w528[52] = |(datain[103:100] ^ 15);
  assign w528[53] = |(datain[99:96] ^ 10);
  assign w528[54] = |(datain[95:92] ^ 12);
  assign w528[55] = |(datain[91:88] ^ 3);
  assign comp[528] = ~(|w528);
  wire [48-1:0] w529;
  assign w529[0] = |(datain[311:308] ^ 14);
  assign w529[1] = |(datain[307:304] ^ 8);
  assign w529[2] = |(datain[303:300] ^ 0);
  assign w529[3] = |(datain[299:296] ^ 0);
  assign w529[4] = |(datain[295:292] ^ 0);
  assign w529[5] = |(datain[291:288] ^ 0);
  assign w529[6] = |(datain[287:284] ^ 5);
  assign w529[7] = |(datain[283:280] ^ 15);
  assign w529[8] = |(datain[279:276] ^ 8);
  assign w529[9] = |(datain[275:272] ^ 1);
  assign w529[10] = |(datain[271:268] ^ 14);
  assign w529[11] = |(datain[267:264] ^ 15);
  assign w529[12] = |(datain[263:260] ^ 0);
  assign w529[13] = |(datain[259:256] ^ 7);
  assign w529[14] = |(datain[255:252] ^ 0);
  assign w529[15] = |(datain[251:248] ^ 1);
  assign w529[16] = |(datain[247:244] ^ 14);
  assign w529[17] = |(datain[243:240] ^ 8);
  assign w529[18] = |(datain[239:236] ^ 0);
  assign w529[19] = |(datain[235:232] ^ 2);
  assign w529[20] = |(datain[231:228] ^ 0);
  assign w529[21] = |(datain[227:224] ^ 0);
  assign w529[22] = |(datain[223:220] ^ 14);
  assign w529[23] = |(datain[219:216] ^ 11);
  assign w529[24] = |(datain[215:212] ^ 1);
  assign w529[25] = |(datain[211:208] ^ 2);
  assign w529[26] = |(datain[207:204] ^ 8);
  assign w529[27] = |(datain[203:200] ^ 13);
  assign w529[28] = |(datain[199:196] ^ 11);
  assign w529[29] = |(datain[195:192] ^ 5);
  assign w529[30] = |(datain[191:188] ^ 2);
  assign w529[31] = |(datain[187:184] ^ 3);
  assign w529[32] = |(datain[183:180] ^ 0);
  assign w529[33] = |(datain[179:176] ^ 1);
  assign w529[34] = |(datain[175:172] ^ 11);
  assign w529[35] = |(datain[171:168] ^ 9);
  assign w529[36] = |(datain[167:164] ^ 11);
  assign w529[37] = |(datain[163:160] ^ 6);
  assign w529[38] = |(datain[159:156] ^ 0);
  assign w529[39] = |(datain[155:152] ^ 3);
  assign w529[40] = |(datain[151:148] ^ 8);
  assign w529[41] = |(datain[147:144] ^ 12);
  assign w529[42] = |(datain[143:140] ^ 12);
  assign w529[43] = |(datain[139:136] ^ 8);
  assign w529[44] = |(datain[135:132] ^ 8);
  assign w529[45] = |(datain[131:128] ^ 14);
  assign w529[46] = |(datain[127:124] ^ 13);
  assign w529[47] = |(datain[123:120] ^ 8);
  assign comp[529] = ~(|w529);
  wire [44-1:0] w530;
  assign w530[0] = |(datain[311:308] ^ 14);
  assign w530[1] = |(datain[307:304] ^ 8);
  assign w530[2] = |(datain[303:300] ^ 0);
  assign w530[3] = |(datain[299:296] ^ 0);
  assign w530[4] = |(datain[295:292] ^ 0);
  assign w530[5] = |(datain[291:288] ^ 0);
  assign w530[6] = |(datain[287:284] ^ 11);
  assign w530[7] = |(datain[283:280] ^ 9);
  assign w530[8] = |(datain[279:276] ^ 1);
  assign w530[9] = |(datain[275:272] ^ 3);
  assign w530[10] = |(datain[271:268] ^ 0);
  assign w530[11] = |(datain[267:264] ^ 1);
  assign w530[12] = |(datain[263:260] ^ 5);
  assign w530[13] = |(datain[259:256] ^ 14);
  assign w530[14] = |(datain[255:252] ^ 8);
  assign w530[15] = |(datain[251:248] ^ 1);
  assign w530[16] = |(datain[247:244] ^ 14);
  assign w530[17] = |(datain[243:240] ^ 14);
  assign w530[18] = |(datain[239:236] ^ 2);
  assign w530[19] = |(datain[235:232] ^ 1);
  assign w530[20] = |(datain[231:228] ^ 0);
  assign w530[21] = |(datain[227:224] ^ 2);
  assign w530[22] = |(datain[223:220] ^ 8);
  assign w530[23] = |(datain[219:216] ^ 13);
  assign w530[24] = |(datain[215:212] ^ 11);
  assign w530[25] = |(datain[211:208] ^ 12);
  assign w530[26] = |(datain[207:204] ^ 0);
  assign w530[27] = |(datain[203:200] ^ 11);
  assign w530[28] = |(datain[199:196] ^ 0);
  assign w530[29] = |(datain[195:192] ^ 1);
  assign w530[30] = |(datain[191:188] ^ 8);
  assign w530[31] = |(datain[187:184] ^ 0);
  assign w530[32] = |(datain[183:180] ^ 3);
  assign w530[33] = |(datain[179:176] ^ 5);
  assign w530[34] = |(datain[175:172] ^ 5);
  assign w530[35] = |(datain[171:168] ^ 1);
  assign w530[36] = |(datain[167:164] ^ 4);
  assign w530[37] = |(datain[163:160] ^ 7);
  assign w530[38] = |(datain[159:156] ^ 14);
  assign w530[39] = |(datain[155:152] ^ 2);
  assign w530[40] = |(datain[151:148] ^ 15);
  assign w530[41] = |(datain[147:144] ^ 10);
  assign w530[42] = |(datain[143:140] ^ 12);
  assign w530[43] = |(datain[139:136] ^ 3);
  assign comp[530] = ~(|w530);
  wire [42-1:0] w531;
  assign w531[0] = |(datain[311:308] ^ 0);
  assign w531[1] = |(datain[307:304] ^ 1);
  assign w531[2] = |(datain[303:300] ^ 8);
  assign w531[3] = |(datain[299:296] ^ 1);
  assign w531[4] = |(datain[295:292] ^ 15);
  assign w531[5] = |(datain[291:288] ^ 12);
  assign w531[6] = |(datain[287:284] ^ 4);
  assign w531[7] = |(datain[283:280] ^ 15);
  assign w531[8] = |(datain[279:276] ^ 5);
  assign w531[9] = |(datain[275:272] ^ 0);
  assign w531[10] = |(datain[271:268] ^ 7);
  assign w531[11] = |(datain[267:264] ^ 4);
  assign w531[12] = |(datain[263:260] ^ 0);
  assign w531[13] = |(datain[259:256] ^ 11);
  assign w531[14] = |(datain[255:252] ^ 8);
  assign w531[15] = |(datain[251:248] ^ 13);
  assign w531[16] = |(datain[247:244] ^ 11);
  assign w531[17] = |(datain[243:240] ^ 6);
  assign w531[18] = |(datain[239:236] ^ 8);
  assign w531[19] = |(datain[235:232] ^ 6);
  assign w531[20] = |(datain[231:228] ^ 0);
  assign w531[21] = |(datain[227:224] ^ 1);
  assign w531[22] = |(datain[223:220] ^ 11);
  assign w531[23] = |(datain[219:216] ^ 15);
  assign w531[24] = |(datain[215:212] ^ 0);
  assign w531[25] = |(datain[211:208] ^ 0);
  assign w531[26] = |(datain[207:204] ^ 0);
  assign w531[27] = |(datain[203:200] ^ 1);
  assign w531[28] = |(datain[199:196] ^ 5);
  assign w531[29] = |(datain[195:192] ^ 7);
  assign w531[30] = |(datain[191:188] ^ 10);
  assign w531[31] = |(datain[187:184] ^ 4);
  assign w531[32] = |(datain[183:180] ^ 14);
  assign w531[33] = |(datain[179:176] ^ 11);
  assign w531[34] = |(datain[175:172] ^ 1);
  assign w531[35] = |(datain[171:168] ^ 1);
  assign w531[36] = |(datain[167:164] ^ 1);
  assign w531[37] = |(datain[163:160] ^ 14);
  assign w531[38] = |(datain[159:156] ^ 0);
  assign w531[39] = |(datain[155:152] ^ 6);
  assign w531[40] = |(datain[151:148] ^ 0);
  assign w531[41] = |(datain[147:144] ^ 14);
  assign comp[531] = ~(|w531);
  wire [54-1:0] w532;
  assign w532[0] = |(datain[311:308] ^ 14);
  assign w532[1] = |(datain[307:304] ^ 8);
  assign w532[2] = |(datain[303:300] ^ 0);
  assign w532[3] = |(datain[299:296] ^ 0);
  assign w532[4] = |(datain[295:292] ^ 0);
  assign w532[5] = |(datain[291:288] ^ 0);
  assign w532[6] = |(datain[287:284] ^ 5);
  assign w532[7] = |(datain[283:280] ^ 13);
  assign w532[8] = |(datain[279:276] ^ 8);
  assign w532[9] = |(datain[275:272] ^ 1);
  assign w532[10] = |(datain[271:268] ^ 14);
  assign w532[11] = |(datain[267:264] ^ 13);
  assign w532[12] = |(datain[263:260] ^ 0);
  assign w532[13] = |(datain[259:256] ^ 6);
  assign w532[14] = |(datain[255:252] ^ 0);
  assign w532[15] = |(datain[251:248] ^ 1);
  assign w532[16] = |(datain[247:244] ^ 8);
  assign w532[17] = |(datain[243:240] ^ 1);
  assign w532[18] = |(datain[239:236] ^ 15);
  assign w532[19] = |(datain[235:232] ^ 12);
  assign w532[20] = |(datain[231:228] ^ 4);
  assign w532[21] = |(datain[227:224] ^ 15);
  assign w532[22] = |(datain[223:220] ^ 5);
  assign w532[23] = |(datain[219:216] ^ 0);
  assign w532[24] = |(datain[215:212] ^ 7);
  assign w532[25] = |(datain[211:208] ^ 4);
  assign w532[26] = |(datain[207:204] ^ 0);
  assign w532[27] = |(datain[203:200] ^ 11);
  assign w532[28] = |(datain[199:196] ^ 8);
  assign w532[29] = |(datain[195:192] ^ 13);
  assign w532[30] = |(datain[191:188] ^ 11);
  assign w532[31] = |(datain[187:184] ^ 6);
  assign w532[32] = |(datain[183:180] ^ 8);
  assign w532[33] = |(datain[179:176] ^ 6);
  assign w532[34] = |(datain[175:172] ^ 0);
  assign w532[35] = |(datain[171:168] ^ 1);
  assign w532[36] = |(datain[167:164] ^ 11);
  assign w532[37] = |(datain[163:160] ^ 15);
  assign w532[38] = |(datain[159:156] ^ 0);
  assign w532[39] = |(datain[155:152] ^ 0);
  assign w532[40] = |(datain[151:148] ^ 0);
  assign w532[41] = |(datain[147:144] ^ 1);
  assign w532[42] = |(datain[143:140] ^ 5);
  assign w532[43] = |(datain[139:136] ^ 7);
  assign w532[44] = |(datain[135:132] ^ 10);
  assign w532[45] = |(datain[131:128] ^ 4);
  assign w532[46] = |(datain[127:124] ^ 14);
  assign w532[47] = |(datain[123:120] ^ 11);
  assign w532[48] = |(datain[119:116] ^ 1);
  assign w532[49] = |(datain[115:112] ^ 1);
  assign w532[50] = |(datain[111:108] ^ 1);
  assign w532[51] = |(datain[107:104] ^ 14);
  assign w532[52] = |(datain[103:100] ^ 0);
  assign w532[53] = |(datain[99:96] ^ 6);
  assign comp[532] = ~(|w532);
  wire [44-1:0] w533;
  assign w533[0] = |(datain[311:308] ^ 0);
  assign w533[1] = |(datain[307:304] ^ 5);
  assign w533[2] = |(datain[303:300] ^ 1);
  assign w533[3] = |(datain[299:296] ^ 0);
  assign w533[4] = |(datain[295:292] ^ 0);
  assign w533[5] = |(datain[291:288] ^ 0);
  assign w533[6] = |(datain[287:284] ^ 3);
  assign w533[7] = |(datain[283:280] ^ 3);
  assign w533[8] = |(datain[279:276] ^ 13);
  assign w533[9] = |(datain[275:272] ^ 11);
  assign w533[10] = |(datain[271:268] ^ 4);
  assign w533[11] = |(datain[267:264] ^ 11);
  assign w533[12] = |(datain[263:260] ^ 8);
  assign w533[13] = |(datain[259:256] ^ 11);
  assign w533[14] = |(datain[255:252] ^ 14);
  assign w533[15] = |(datain[251:248] ^ 3);
  assign w533[16] = |(datain[247:244] ^ 8);
  assign w533[17] = |(datain[243:240] ^ 14);
  assign w533[18] = |(datain[239:236] ^ 13);
  assign w533[19] = |(datain[235:232] ^ 0);
  assign w533[20] = |(datain[231:228] ^ 14);
  assign w533[21] = |(datain[227:224] ^ 8);
  assign w533[22] = |(datain[223:220] ^ 0);
  assign w533[23] = |(datain[219:216] ^ 5);
  assign w533[24] = |(datain[215:212] ^ 0);
  assign w533[25] = |(datain[211:208] ^ 2);
  assign w533[26] = |(datain[207:204] ^ 10);
  assign w533[27] = |(datain[203:200] ^ 1);
  assign w533[28] = |(datain[199:196] ^ 15);
  assign w533[29] = |(datain[195:192] ^ 11);
  assign w533[30] = |(datain[191:188] ^ 0);
  assign w533[31] = |(datain[187:184] ^ 2);
  assign w533[32] = |(datain[183:180] ^ 8);
  assign w533[33] = |(datain[179:176] ^ 12);
  assign w533[34] = |(datain[175:172] ^ 12);
  assign w533[35] = |(datain[171:168] ^ 3);
  assign w533[36] = |(datain[167:164] ^ 0);
  assign w533[37] = |(datain[163:160] ^ 3);
  assign w533[38] = |(datain[159:156] ^ 12);
  assign w533[39] = |(datain[155:152] ^ 3);
  assign w533[40] = |(datain[151:148] ^ 10);
  assign w533[41] = |(datain[147:144] ^ 3);
  assign w533[42] = |(datain[143:140] ^ 5);
  assign w533[43] = |(datain[139:136] ^ 4);
  assign comp[533] = ~(|w533);
  wire [42-1:0] w534;
  assign w534[0] = |(datain[311:308] ^ 0);
  assign w534[1] = |(datain[307:304] ^ 6);
  assign w534[2] = |(datain[303:300] ^ 7);
  assign w534[3] = |(datain[299:296] ^ 4);
  assign w534[4] = |(datain[295:292] ^ 0);
  assign w534[5] = |(datain[291:288] ^ 3);
  assign w534[6] = |(datain[287:284] ^ 8);
  assign w534[7] = |(datain[283:280] ^ 12);
  assign w534[8] = |(datain[279:276] ^ 1);
  assign w534[9] = |(datain[275:272] ^ 6);
  assign w534[10] = |(datain[271:268] ^ 7);
  assign w534[11] = |(datain[267:264] ^ 6);
  assign w534[12] = |(datain[263:260] ^ 0);
  assign w534[13] = |(datain[259:256] ^ 3);
  assign w534[14] = |(datain[255:252] ^ 8);
  assign w534[15] = |(datain[251:248] ^ 9);
  assign w534[16] = |(datain[247:244] ^ 2);
  assign w534[17] = |(datain[243:240] ^ 6);
  assign w534[18] = |(datain[239:236] ^ 7);
  assign w534[19] = |(datain[235:232] ^ 8);
  assign w534[20] = |(datain[231:228] ^ 0);
  assign w534[21] = |(datain[227:224] ^ 3);
  assign w534[22] = |(datain[223:220] ^ 8);
  assign w534[23] = |(datain[219:216] ^ 12);
  assign w534[24] = |(datain[215:212] ^ 12);
  assign w534[25] = |(datain[211:208] ^ 8);
  assign w534[26] = |(datain[207:204] ^ 0);
  assign w534[27] = |(datain[203:200] ^ 5);
  assign w534[28] = |(datain[199:196] ^ 1);
  assign w534[29] = |(datain[195:192] ^ 0);
  assign w534[30] = |(datain[191:188] ^ 0);
  assign w534[31] = |(datain[187:184] ^ 0);
  assign w534[32] = |(datain[183:180] ^ 3);
  assign w534[33] = |(datain[179:176] ^ 3);
  assign w534[34] = |(datain[175:172] ^ 13);
  assign w534[35] = |(datain[171:168] ^ 11);
  assign w534[36] = |(datain[167:164] ^ 4);
  assign w534[37] = |(datain[163:160] ^ 11);
  assign w534[38] = |(datain[159:156] ^ 8);
  assign w534[39] = |(datain[155:152] ^ 11);
  assign w534[40] = |(datain[151:148] ^ 14);
  assign w534[41] = |(datain[147:144] ^ 3);
  assign comp[534] = ~(|w534);
  wire [28-1:0] w535;
  assign w535[0] = |(datain[311:308] ^ 1);
  assign w535[1] = |(datain[307:304] ^ 2);
  assign w535[2] = |(datain[303:300] ^ 0);
  assign w535[3] = |(datain[299:296] ^ 1);
  assign w535[4] = |(datain[295:292] ^ 11);
  assign w535[5] = |(datain[291:288] ^ 15);
  assign w535[6] = |(datain[287:284] ^ 1);
  assign w535[7] = |(datain[283:280] ^ 10);
  assign w535[8] = |(datain[279:276] ^ 15);
  assign w535[9] = |(datain[275:272] ^ 15);
  assign w535[10] = |(datain[271:268] ^ 8);
  assign w535[11] = |(datain[267:264] ^ 1);
  assign w535[12] = |(datain[263:260] ^ 3);
  assign w535[13] = |(datain[259:256] ^ 4);
  assign w535[14] = |(datain[255:252] ^ 0);
  assign w535[15] = |(datain[251:248] ^ 0);
  assign w535[16] = |(datain[247:244] ^ 0);
  assign w535[17] = |(datain[243:240] ^ 0);
  assign w535[18] = |(datain[239:236] ^ 4);
  assign w535[19] = |(datain[235:232] ^ 6);
  assign w535[20] = |(datain[231:228] ^ 4);
  assign w535[21] = |(datain[227:224] ^ 6);
  assign w535[22] = |(datain[223:220] ^ 4);
  assign w535[23] = |(datain[219:216] ^ 7);
  assign w535[24] = |(datain[215:212] ^ 7);
  assign w535[25] = |(datain[211:208] ^ 5);
  assign w535[26] = |(datain[207:204] ^ 15);
  assign w535[27] = |(datain[203:200] ^ 7);
  assign comp[535] = ~(|w535);
  wire [34-1:0] w536;
  assign w536[0] = |(datain[311:308] ^ 1);
  assign w536[1] = |(datain[307:304] ^ 7);
  assign w536[2] = |(datain[303:300] ^ 0);
  assign w536[3] = |(datain[299:296] ^ 1);
  assign w536[4] = |(datain[295:292] ^ 11);
  assign w536[5] = |(datain[291:288] ^ 13);
  assign w536[6] = |(datain[287:284] ^ 8);
  assign w536[7] = |(datain[283:280] ^ 9);
  assign w536[8] = |(datain[279:276] ^ 15);
  assign w536[9] = |(datain[275:272] ^ 14);
  assign w536[10] = |(datain[271:268] ^ 14);
  assign w536[11] = |(datain[267:264] ^ 2);
  assign w536[12] = |(datain[263:260] ^ 15);
  assign w536[13] = |(datain[259:256] ^ 14);
  assign w536[14] = |(datain[255:252] ^ 2);
  assign w536[15] = |(datain[251:248] ^ 14);
  assign w536[16] = |(datain[247:244] ^ 8);
  assign w536[17] = |(datain[243:240] ^ 1);
  assign w536[18] = |(datain[239:236] ^ 2);
  assign w536[19] = |(datain[235:232] ^ 12);
  assign w536[20] = |(datain[231:228] ^ 0);
  assign w536[21] = |(datain[227:224] ^ 0);
  assign w536[22] = |(datain[223:220] ^ 0);
  assign w536[23] = |(datain[219:216] ^ 0);
  assign w536[24] = |(datain[215:212] ^ 4);
  assign w536[25] = |(datain[211:208] ^ 6);
  assign w536[26] = |(datain[207:204] ^ 4);
  assign w536[27] = |(datain[203:200] ^ 6);
  assign w536[28] = |(datain[199:196] ^ 4);
  assign w536[29] = |(datain[195:192] ^ 5);
  assign w536[30] = |(datain[191:188] ^ 7);
  assign w536[31] = |(datain[187:184] ^ 5);
  assign w536[32] = |(datain[183:180] ^ 15);
  assign w536[33] = |(datain[179:176] ^ 6);
  assign comp[536] = ~(|w536);
  wire [32-1:0] w537;
  assign w537[0] = |(datain[311:308] ^ 15);
  assign w537[1] = |(datain[307:304] ^ 10);
  assign w537[2] = |(datain[303:300] ^ 15);
  assign w537[3] = |(datain[299:296] ^ 14);
  assign w537[4] = |(datain[295:292] ^ 11);
  assign w537[5] = |(datain[291:288] ^ 13);
  assign w537[6] = |(datain[287:284] ^ 1);
  assign w537[7] = |(datain[283:280] ^ 1);
  assign w537[8] = |(datain[279:276] ^ 0);
  assign w537[9] = |(datain[275:272] ^ 1);
  assign w537[10] = |(datain[271:268] ^ 2);
  assign w537[11] = |(datain[267:264] ^ 14);
  assign w537[12] = |(datain[263:260] ^ 8);
  assign w537[13] = |(datain[259:256] ^ 1);
  assign w537[14] = |(datain[255:252] ^ 7);
  assign w537[15] = |(datain[251:248] ^ 6);
  assign w537[16] = |(datain[247:244] ^ 0);
  assign w537[17] = |(datain[243:240] ^ 0);
  assign w537[18] = |(datain[239:236] ^ 0);
  assign w537[19] = |(datain[235:232] ^ 0);
  assign w537[20] = |(datain[231:228] ^ 0);
  assign w537[21] = |(datain[227:224] ^ 0);
  assign w537[22] = |(datain[223:220] ^ 4);
  assign w537[23] = |(datain[219:216] ^ 5);
  assign w537[24] = |(datain[215:212] ^ 4);
  assign w537[25] = |(datain[211:208] ^ 5);
  assign w537[26] = |(datain[207:204] ^ 4);
  assign w537[27] = |(datain[203:200] ^ 2);
  assign w537[28] = |(datain[199:196] ^ 7);
  assign w537[29] = |(datain[195:192] ^ 5);
  assign w537[30] = |(datain[191:188] ^ 15);
  assign w537[31] = |(datain[187:184] ^ 5);
  assign comp[537] = ~(|w537);
  wire [46-1:0] w538;
  assign w538[0] = |(datain[311:308] ^ 14);
  assign w538[1] = |(datain[307:304] ^ 8);
  assign w538[2] = |(datain[303:300] ^ 0);
  assign w538[3] = |(datain[299:296] ^ 0);
  assign w538[4] = |(datain[295:292] ^ 0);
  assign w538[5] = |(datain[291:288] ^ 0);
  assign w538[6] = |(datain[287:284] ^ 5);
  assign w538[7] = |(datain[283:280] ^ 8);
  assign w538[8] = |(datain[279:276] ^ 9);
  assign w538[9] = |(datain[275:272] ^ 6);
  assign w538[10] = |(datain[271:268] ^ 8);
  assign w538[11] = |(datain[267:264] ^ 1);
  assign w538[12] = |(datain[263:260] ^ 14);
  assign w538[13] = |(datain[259:256] ^ 14);
  assign w538[14] = |(datain[255:252] ^ 1);
  assign w538[15] = |(datain[251:248] ^ 9);
  assign w538[16] = |(datain[247:244] ^ 0);
  assign w538[17] = |(datain[243:240] ^ 1);
  assign w538[18] = |(datain[239:236] ^ 8);
  assign w538[19] = |(datain[235:232] ^ 13);
  assign w538[20] = |(datain[231:228] ^ 11);
  assign w538[21] = |(datain[227:224] ^ 12);
  assign w538[22] = |(datain[223:220] ^ 2);
  assign w538[23] = |(datain[219:216] ^ 13);
  assign w538[24] = |(datain[215:212] ^ 0);
  assign w538[25] = |(datain[211:208] ^ 1);
  assign w538[26] = |(datain[207:204] ^ 11);
  assign w538[27] = |(datain[203:200] ^ 9);
  assign w538[28] = |(datain[199:196] ^ 13);
  assign w538[29] = |(datain[195:192] ^ 10);
  assign w538[30] = |(datain[191:188] ^ 0);
  assign w538[31] = |(datain[187:184] ^ 2);
  assign w538[32] = |(datain[183:180] ^ 8);
  assign w538[33] = |(datain[179:176] ^ 0);
  assign w538[34] = |(datain[175:172] ^ 3);
  assign w538[35] = |(datain[171:168] ^ 5);
  assign w538[36] = |(datain[167:164] ^ 0);
  assign w538[37] = |(datain[163:160] ^ 1);
  assign w538[38] = |(datain[159:156] ^ 4);
  assign w538[39] = |(datain[155:152] ^ 7);
  assign w538[40] = |(datain[151:148] ^ 14);
  assign w538[41] = |(datain[147:144] ^ 2);
  assign w538[42] = |(datain[143:140] ^ 15);
  assign w538[43] = |(datain[139:136] ^ 10);
  assign w538[44] = |(datain[135:132] ^ 12);
  assign w538[45] = |(datain[131:128] ^ 3);
  assign comp[538] = ~(|w538);
  wire [36-1:0] w539;
  assign w539[0] = |(datain[311:308] ^ 11);
  assign w539[1] = |(datain[307:304] ^ 10);
  assign w539[2] = |(datain[303:300] ^ 6);
  assign w539[3] = |(datain[299:296] ^ 12);
  assign w539[4] = |(datain[295:292] ^ 15);
  assign w539[5] = |(datain[291:288] ^ 14);
  assign w539[6] = |(datain[287:284] ^ 11);
  assign w539[7] = |(datain[283:280] ^ 15);
  assign w539[8] = |(datain[279:276] ^ 1);
  assign w539[9] = |(datain[275:272] ^ 1);
  assign w539[10] = |(datain[271:268] ^ 0);
  assign w539[11] = |(datain[267:264] ^ 0);
  assign w539[12] = |(datain[263:260] ^ 14);
  assign w539[13] = |(datain[259:256] ^ 2);
  assign w539[14] = |(datain[255:252] ^ 15);
  assign w539[15] = |(datain[251:248] ^ 14);
  assign w539[16] = |(datain[247:244] ^ 4);
  assign w539[17] = |(datain[243:240] ^ 7);
  assign w539[18] = |(datain[239:236] ^ 2);
  assign w539[19] = |(datain[235:232] ^ 14);
  assign w539[20] = |(datain[231:228] ^ 8);
  assign w539[21] = |(datain[227:224] ^ 1);
  assign w539[22] = |(datain[223:220] ^ 0);
  assign w539[23] = |(datain[219:216] ^ 5);
  assign w539[24] = |(datain[215:212] ^ 0);
  assign w539[25] = |(datain[211:208] ^ 0);
  assign w539[26] = |(datain[207:204] ^ 0);
  assign w539[27] = |(datain[203:200] ^ 0);
  assign w539[28] = |(datain[199:196] ^ 4);
  assign w539[29] = |(datain[195:192] ^ 7);
  assign w539[30] = |(datain[191:188] ^ 4);
  assign w539[31] = |(datain[187:184] ^ 2);
  assign w539[32] = |(datain[183:180] ^ 7);
  assign w539[33] = |(datain[179:176] ^ 5);
  assign w539[34] = |(datain[175:172] ^ 15);
  assign w539[35] = |(datain[171:168] ^ 6);
  assign comp[539] = ~(|w539);
  wire [40-1:0] w540;
  assign w540[0] = |(datain[311:308] ^ 7);
  assign w540[1] = |(datain[307:304] ^ 9);
  assign w540[2] = |(datain[303:300] ^ 7);
  assign w540[3] = |(datain[299:296] ^ 10);
  assign w540[4] = |(datain[295:292] ^ 12);
  assign w540[5] = |(datain[291:288] ^ 13);
  assign w540[6] = |(datain[287:284] ^ 2);
  assign w540[7] = |(datain[283:280] ^ 1);
  assign w540[8] = |(datain[279:276] ^ 3);
  assign w540[9] = |(datain[275:272] ^ 13);
  assign w540[10] = |(datain[271:268] ^ 5);
  assign w540[11] = |(datain[267:264] ^ 9);
  assign w540[12] = |(datain[263:260] ^ 5);
  assign w540[13] = |(datain[259:256] ^ 10);
  assign w540[14] = |(datain[255:252] ^ 7);
  assign w540[15] = |(datain[251:248] ^ 4);
  assign w540[16] = |(datain[247:244] ^ 5);
  assign w540[17] = |(datain[243:240] ^ 8);
  assign w540[18] = |(datain[239:236] ^ 3);
  assign w540[19] = |(datain[235:232] ^ 3);
  assign w540[20] = |(datain[231:228] ^ 12);
  assign w540[21] = |(datain[227:224] ^ 0);
  assign w540[22] = |(datain[223:220] ^ 8);
  assign w540[23] = |(datain[219:216] ^ 14);
  assign w540[24] = |(datain[215:212] ^ 13);
  assign w540[25] = |(datain[211:208] ^ 8);
  assign w540[26] = |(datain[207:204] ^ 8);
  assign w540[27] = |(datain[203:200] ^ 12);
  assign w540[28] = |(datain[199:196] ^ 12);
  assign w540[29] = |(datain[195:192] ^ 0);
  assign w540[30] = |(datain[191:188] ^ 4);
  assign w540[31] = |(datain[187:184] ^ 8);
  assign w540[32] = |(datain[183:180] ^ 8);
  assign w540[33] = |(datain[179:176] ^ 14);
  assign w540[34] = |(datain[175:172] ^ 12);
  assign w540[35] = |(datain[171:168] ^ 0);
  assign w540[36] = |(datain[167:164] ^ 10);
  assign w540[37] = |(datain[163:160] ^ 1);
  assign w540[38] = |(datain[159:156] ^ 8);
  assign w540[39] = |(datain[155:152] ^ 4);
  assign comp[540] = ~(|w540);
  wire [46-1:0] w541;
  assign w541[0] = |(datain[311:308] ^ 5);
  assign w541[1] = |(datain[307:304] ^ 1);
  assign w541[2] = |(datain[303:300] ^ 5);
  assign w541[3] = |(datain[299:296] ^ 2);
  assign w541[4] = |(datain[295:292] ^ 5);
  assign w541[5] = |(datain[291:288] ^ 0);
  assign w541[6] = |(datain[287:284] ^ 14);
  assign w541[7] = |(datain[283:280] ^ 8);
  assign w541[8] = |(datain[279:276] ^ 6);
  assign w541[9] = |(datain[275:272] ^ 13);
  assign w541[10] = |(datain[271:268] ^ 15);
  assign w541[11] = |(datain[267:264] ^ 13);
  assign w541[12] = |(datain[263:260] ^ 2);
  assign w541[13] = |(datain[259:256] ^ 14);
  assign w541[14] = |(datain[255:252] ^ 8);
  assign w541[15] = |(datain[251:248] ^ 3);
  assign w541[16] = |(datain[247:244] ^ 8);
  assign w541[17] = |(datain[243:240] ^ 4);
  assign w541[18] = |(datain[239:236] ^ 12);
  assign w541[19] = |(datain[235:232] ^ 3);
  assign w541[20] = |(datain[231:228] ^ 0);
  assign w541[21] = |(datain[227:224] ^ 3);
  assign w541[22] = |(datain[223:220] ^ 0);
  assign w541[23] = |(datain[219:216] ^ 1);
  assign w541[24] = |(datain[215:212] ^ 14);
  assign w541[25] = |(datain[211:208] ^ 8);
  assign w541[26] = |(datain[207:204] ^ 2);
  assign w541[27] = |(datain[203:200] ^ 2);
  assign w541[28] = |(datain[199:196] ^ 15);
  assign w541[29] = |(datain[195:192] ^ 15);
  assign w541[30] = |(datain[191:188] ^ 14);
  assign w541[31] = |(datain[187:184] ^ 8);
  assign w541[32] = |(datain[183:180] ^ 13);
  assign w541[33] = |(datain[179:176] ^ 8);
  assign w541[34] = |(datain[175:172] ^ 15);
  assign w541[35] = |(datain[171:168] ^ 15);
  assign w541[36] = |(datain[167:164] ^ 5);
  assign w541[37] = |(datain[163:160] ^ 8);
  assign w541[38] = |(datain[159:156] ^ 5);
  assign w541[39] = |(datain[155:152] ^ 10);
  assign w541[40] = |(datain[151:148] ^ 5);
  assign w541[41] = |(datain[147:144] ^ 9);
  assign w541[42] = |(datain[143:140] ^ 5);
  assign w541[43] = |(datain[139:136] ^ 11);
  assign w541[44] = |(datain[135:132] ^ 12);
  assign w541[45] = |(datain[131:128] ^ 13);
  assign comp[541] = ~(|w541);
  wire [46-1:0] w542;
  assign w542[0] = |(datain[311:308] ^ 4);
  assign w542[1] = |(datain[307:304] ^ 0);
  assign w542[2] = |(datain[303:300] ^ 8);
  assign w542[3] = |(datain[299:296] ^ 11);
  assign w542[4] = |(datain[295:292] ^ 9);
  assign w542[5] = |(datain[291:288] ^ 12);
  assign w542[6] = |(datain[287:284] ^ 3);
  assign w542[7] = |(datain[283:280] ^ 0);
  assign w542[8] = |(datain[279:276] ^ 0);
  assign w542[9] = |(datain[275:272] ^ 4);
  assign w542[10] = |(datain[271:268] ^ 11);
  assign w542[11] = |(datain[267:264] ^ 9);
  assign w542[12] = |(datain[263:260] ^ 14);
  assign w542[13] = |(datain[259:256] ^ 1);
  assign w542[14] = |(datain[255:252] ^ 0);
  assign w542[15] = |(datain[251:248] ^ 2);
  assign w542[16] = |(datain[247:244] ^ 8);
  assign w542[17] = |(datain[243:240] ^ 13);
  assign w542[18] = |(datain[239:236] ^ 9);
  assign w542[19] = |(datain[235:232] ^ 4);
  assign w542[20] = |(datain[231:228] ^ 0);
  assign w542[21] = |(datain[227:224] ^ 14);
  assign w542[22] = |(datain[223:220] ^ 0);
  assign w542[23] = |(datain[219:216] ^ 1);
  assign w542[24] = |(datain[215:212] ^ 12);
  assign w542[25] = |(datain[211:208] ^ 13);
  assign w542[26] = |(datain[207:204] ^ 2);
  assign w542[27] = |(datain[203:200] ^ 1);
  assign w542[28] = |(datain[199:196] ^ 14);
  assign w542[29] = |(datain[195:192] ^ 8);
  assign w542[30] = |(datain[191:188] ^ 13);
  assign w542[31] = |(datain[187:184] ^ 6);
  assign w542[32] = |(datain[183:180] ^ 15);
  assign w542[33] = |(datain[179:176] ^ 15);
  assign w542[34] = |(datain[175:172] ^ 14);
  assign w542[35] = |(datain[171:168] ^ 8);
  assign w542[36] = |(datain[167:164] ^ 12);
  assign w542[37] = |(datain[163:160] ^ 3);
  assign w542[38] = |(datain[159:156] ^ 15);
  assign w542[39] = |(datain[155:152] ^ 15);
  assign w542[40] = |(datain[151:148] ^ 12);
  assign w542[41] = |(datain[147:144] ^ 3);
  assign w542[42] = |(datain[143:140] ^ 4);
  assign w542[43] = |(datain[139:136] ^ 9);
  assign w542[44] = |(datain[135:132] ^ 6);
  assign w542[45] = |(datain[131:128] ^ 13);
  assign comp[542] = ~(|w542);
  wire [60-1:0] w543;
  assign w543[0] = |(datain[311:308] ^ 8);
  assign w543[1] = |(datain[307:304] ^ 14);
  assign w543[2] = |(datain[303:300] ^ 11);
  assign w543[3] = |(datain[299:296] ^ 15);
  assign w543[4] = |(datain[295:292] ^ 1);
  assign w543[5] = |(datain[291:288] ^ 14);
  assign w543[6] = |(datain[287:284] ^ 0);
  assign w543[7] = |(datain[283:280] ^ 2);
  assign w543[8] = |(datain[279:276] ^ 11);
  assign w543[9] = |(datain[275:272] ^ 10);
  assign w543[10] = |(datain[271:268] ^ 9);
  assign w543[11] = |(datain[267:264] ^ 0);
  assign w543[12] = |(datain[263:260] ^ 0);
  assign w543[13] = |(datain[259:256] ^ 1);
  assign w543[14] = |(datain[255:252] ^ 8);
  assign w543[15] = |(datain[251:248] ^ 9);
  assign w543[16] = |(datain[247:244] ^ 0);
  assign w543[17] = |(datain[243:240] ^ 6);
  assign w543[18] = |(datain[239:236] ^ 12);
  assign w543[19] = |(datain[235:232] ^ 3);
  assign w543[20] = |(datain[231:228] ^ 12);
  assign w543[21] = |(datain[227:224] ^ 3);
  assign w543[22] = |(datain[223:220] ^ 0);
  assign w543[23] = |(datain[219:216] ^ 7);
  assign w543[24] = |(datain[215:212] ^ 10);
  assign w543[25] = |(datain[211:208] ^ 9);
  assign w543[26] = |(datain[207:204] ^ 14);
  assign w543[27] = |(datain[203:200] ^ 1);
  assign w543[28] = |(datain[199:196] ^ 15);
  assign w543[29] = |(datain[195:192] ^ 11);
  assign w543[30] = |(datain[191:188] ^ 12);
  assign w543[31] = |(datain[187:184] ^ 0);
  assign w543[32] = |(datain[183:180] ^ 8);
  assign w543[33] = |(datain[179:176] ^ 13);
  assign w543[34] = |(datain[175:172] ^ 11);
  assign w543[35] = |(datain[171:168] ^ 12);
  assign w543[36] = |(datain[167:164] ^ 1);
  assign w543[37] = |(datain[163:160] ^ 13);
  assign w543[38] = |(datain[159:156] ^ 0);
  assign w543[39] = |(datain[155:152] ^ 1);
  assign w543[40] = |(datain[151:148] ^ 11);
  assign w543[41] = |(datain[147:144] ^ 9);
  assign w543[42] = |(datain[143:140] ^ 10);
  assign w543[43] = |(datain[139:136] ^ 3);
  assign w543[44] = |(datain[135:132] ^ 0);
  assign w543[45] = |(datain[131:128] ^ 2);
  assign w543[46] = |(datain[127:124] ^ 8);
  assign w543[47] = |(datain[123:120] ^ 0);
  assign w543[48] = |(datain[119:116] ^ 3);
  assign w543[49] = |(datain[115:112] ^ 5);
  assign w543[50] = |(datain[111:108] ^ 0);
  assign w543[51] = |(datain[107:104] ^ 3);
  assign w543[52] = |(datain[103:100] ^ 4);
  assign w543[53] = |(datain[99:96] ^ 7);
  assign w543[54] = |(datain[95:92] ^ 14);
  assign w543[55] = |(datain[91:88] ^ 2);
  assign w543[56] = |(datain[87:84] ^ 15);
  assign w543[57] = |(datain[83:80] ^ 10);
  assign w543[58] = |(datain[79:76] ^ 12);
  assign w543[59] = |(datain[75:72] ^ 3);
  assign comp[543] = ~(|w543);
  wire [42-1:0] w544;
  assign w544[0] = |(datain[311:308] ^ 4);
  assign w544[1] = |(datain[307:304] ^ 0);
  assign w544[2] = |(datain[303:300] ^ 8);
  assign w544[3] = |(datain[299:296] ^ 11);
  assign w544[4] = |(datain[295:292] ^ 9);
  assign w544[5] = |(datain[291:288] ^ 12);
  assign w544[6] = |(datain[287:284] ^ 3);
  assign w544[7] = |(datain[283:280] ^ 5);
  assign w544[8] = |(datain[279:276] ^ 0);
  assign w544[9] = |(datain[275:272] ^ 4);
  assign w544[10] = |(datain[271:268] ^ 11);
  assign w544[11] = |(datain[267:264] ^ 9);
  assign w544[12] = |(datain[263:260] ^ 14);
  assign w544[13] = |(datain[259:256] ^ 6);
  assign w544[14] = |(datain[255:252] ^ 0);
  assign w544[15] = |(datain[251:248] ^ 2);
  assign w544[16] = |(datain[247:244] ^ 8);
  assign w544[17] = |(datain[243:240] ^ 13);
  assign w544[18] = |(datain[239:236] ^ 9);
  assign w544[19] = |(datain[235:232] ^ 4);
  assign w544[20] = |(datain[231:228] ^ 0);
  assign w544[21] = |(datain[227:224] ^ 14);
  assign w544[22] = |(datain[223:220] ^ 0);
  assign w544[23] = |(datain[219:216] ^ 1);
  assign w544[24] = |(datain[215:212] ^ 12);
  assign w544[25] = |(datain[211:208] ^ 13);
  assign w544[26] = |(datain[207:204] ^ 2);
  assign w544[27] = |(datain[203:200] ^ 1);
  assign w544[28] = |(datain[199:196] ^ 14);
  assign w544[29] = |(datain[195:192] ^ 8);
  assign w544[30] = |(datain[191:188] ^ 13);
  assign w544[31] = |(datain[187:184] ^ 6);
  assign w544[32] = |(datain[183:180] ^ 15);
  assign w544[33] = |(datain[179:176] ^ 15);
  assign w544[34] = |(datain[175:172] ^ 14);
  assign w544[35] = |(datain[171:168] ^ 8);
  assign w544[36] = |(datain[167:164] ^ 11);
  assign w544[37] = |(datain[163:160] ^ 14);
  assign w544[38] = |(datain[159:156] ^ 15);
  assign w544[39] = |(datain[155:152] ^ 15);
  assign w544[40] = |(datain[151:148] ^ 12);
  assign w544[41] = |(datain[147:144] ^ 3);
  assign comp[544] = ~(|w544);
  wire [50-1:0] w545;
  assign w545[0] = |(datain[311:308] ^ 5);
  assign w545[1] = |(datain[307:304] ^ 14);
  assign w545[2] = |(datain[303:300] ^ 8);
  assign w545[3] = |(datain[299:296] ^ 1);
  assign w545[4] = |(datain[295:292] ^ 14);
  assign w545[5] = |(datain[291:288] ^ 14);
  assign w545[6] = |(datain[287:284] ^ 0);
  assign w545[7] = |(datain[283:280] ^ 6);
  assign w545[8] = |(datain[279:276] ^ 0);
  assign w545[9] = |(datain[275:272] ^ 0);
  assign w545[10] = |(datain[271:268] ^ 8);
  assign w545[11] = |(datain[267:264] ^ 13);
  assign w545[12] = |(datain[263:260] ^ 8);
  assign w545[13] = |(datain[259:256] ^ 4);
  assign w545[14] = |(datain[255:252] ^ 1);
  assign w545[15] = |(datain[251:248] ^ 15);
  assign w545[16] = |(datain[247:244] ^ 0);
  assign w545[17] = |(datain[243:240] ^ 0);
  assign w545[18] = |(datain[239:236] ^ 5);
  assign w545[19] = |(datain[235:232] ^ 0);
  assign w545[20] = |(datain[231:228] ^ 8);
  assign w545[21] = |(datain[227:224] ^ 13);
  assign w545[22] = |(datain[223:220] ^ 11);
  assign w545[23] = |(datain[219:216] ^ 12);
  assign w545[24] = |(datain[215:212] ^ 1);
  assign w545[25] = |(datain[211:208] ^ 15);
  assign w545[26] = |(datain[207:204] ^ 0);
  assign w545[27] = |(datain[203:200] ^ 0);
  assign w545[28] = |(datain[199:196] ^ 11);
  assign w545[29] = |(datain[195:192] ^ 9);
  assign w545[30] = |(datain[191:188] ^ 4);
  assign w545[31] = |(datain[187:184] ^ 12);
  assign w545[32] = |(datain[183:180] ^ 0);
  assign w545[33] = |(datain[179:176] ^ 4);
  assign w545[34] = |(datain[175:172] ^ 2);
  assign w545[35] = |(datain[171:168] ^ 14);
  assign w545[36] = |(datain[167:164] ^ 8);
  assign w545[37] = |(datain[163:160] ^ 0);
  assign w545[38] = |(datain[159:156] ^ 2);
  assign w545[39] = |(datain[155:152] ^ 13);
  assign w545[40] = |(datain[151:148] ^ 2);
  assign w545[41] = |(datain[147:144] ^ 1);
  assign w545[42] = |(datain[143:140] ^ 4);
  assign w545[43] = |(datain[139:136] ^ 7);
  assign w545[44] = |(datain[135:132] ^ 14);
  assign w545[45] = |(datain[131:128] ^ 2);
  assign w545[46] = |(datain[127:124] ^ 15);
  assign w545[47] = |(datain[123:120] ^ 9);
  assign w545[48] = |(datain[119:116] ^ 12);
  assign w545[49] = |(datain[115:112] ^ 3);
  assign comp[545] = ~(|w545);
  wire [44-1:0] w546;
  assign w546[0] = |(datain[311:308] ^ 1);
  assign w546[1] = |(datain[307:304] ^ 5);
  assign w546[2] = |(datain[303:300] ^ 4);
  assign w546[3] = |(datain[299:296] ^ 7);
  assign w546[4] = |(datain[295:292] ^ 14);
  assign w546[5] = |(datain[291:288] ^ 2);
  assign w546[6] = |(datain[287:284] ^ 15);
  assign w546[7] = |(datain[283:280] ^ 10);
  assign w546[8] = |(datain[279:276] ^ 12);
  assign w546[9] = |(datain[275:272] ^ 3);
  assign w546[10] = |(datain[271:268] ^ 9);
  assign w546[11] = |(datain[267:264] ^ 0);
  assign w546[12] = |(datain[263:260] ^ 5);
  assign w546[13] = |(datain[259:256] ^ 0);
  assign w546[14] = |(datain[255:252] ^ 5);
  assign w546[15] = |(datain[251:248] ^ 3);
  assign w546[16] = |(datain[247:244] ^ 5);
  assign w546[17] = |(datain[243:240] ^ 1);
  assign w546[18] = |(datain[239:236] ^ 5);
  assign w546[19] = |(datain[235:232] ^ 2);
  assign w546[20] = |(datain[231:228] ^ 2);
  assign w546[21] = |(datain[227:224] ^ 14);
  assign w546[22] = |(datain[223:220] ^ 8);
  assign w546[23] = |(datain[219:216] ^ 0);
  assign w546[24] = |(datain[215:212] ^ 8);
  assign w546[25] = |(datain[211:208] ^ 4);
  assign w546[26] = |(datain[207:204] ^ 7);
  assign w546[27] = |(datain[203:200] ^ 14);
  assign w546[28] = |(datain[199:196] ^ 0);
  assign w546[29] = |(datain[195:192] ^ 3);
  assign w546[30] = |(datain[191:188] ^ 0);
  assign w546[31] = |(datain[187:184] ^ 2);
  assign w546[32] = |(datain[183:180] ^ 14);
  assign w546[33] = |(datain[179:176] ^ 8);
  assign w546[34] = |(datain[175:172] ^ 6);
  assign w546[35] = |(datain[171:168] ^ 14);
  assign w546[36] = |(datain[167:164] ^ 15);
  assign w546[37] = |(datain[163:160] ^ 15);
  assign w546[38] = |(datain[159:156] ^ 14);
  assign w546[39] = |(datain[155:152] ^ 8);
  assign w546[40] = |(datain[151:148] ^ 13);
  assign w546[41] = |(datain[147:144] ^ 14);
  assign w546[42] = |(datain[143:140] ^ 15);
  assign w546[43] = |(datain[139:136] ^ 15);
  assign comp[546] = ~(|w546);
  wire [34-1:0] w547;
  assign w547[0] = |(datain[311:308] ^ 10);
  assign w547[1] = |(datain[307:304] ^ 6);
  assign w547[2] = |(datain[303:300] ^ 15);
  assign w547[3] = |(datain[299:296] ^ 14);
  assign w547[4] = |(datain[295:292] ^ 14);
  assign w547[5] = |(datain[291:288] ^ 2);
  assign w547[6] = |(datain[287:284] ^ 15);
  assign w547[7] = |(datain[283:280] ^ 14);
  assign w547[8] = |(datain[279:276] ^ 11);
  assign w547[9] = |(datain[275:272] ^ 14);
  assign w547[10] = |(datain[271:268] ^ 1);
  assign w547[11] = |(datain[267:264] ^ 13);
  assign w547[12] = |(datain[263:260] ^ 0);
  assign w547[13] = |(datain[259:256] ^ 0);
  assign w547[14] = |(datain[255:252] ^ 4);
  assign w547[15] = |(datain[251:248] ^ 6);
  assign w547[16] = |(datain[247:244] ^ 2);
  assign w547[17] = |(datain[243:240] ^ 14);
  assign w547[18] = |(datain[239:236] ^ 8);
  assign w547[19] = |(datain[235:232] ^ 1);
  assign w547[20] = |(datain[231:228] ^ 3);
  assign w547[21] = |(datain[227:224] ^ 4);
  assign w547[22] = |(datain[223:220] ^ 8);
  assign w547[23] = |(datain[219:216] ^ 4);
  assign w547[24] = |(datain[215:212] ^ 11);
  assign w547[25] = |(datain[211:208] ^ 14);
  assign w547[26] = |(datain[207:204] ^ 4);
  assign w547[27] = |(datain[203:200] ^ 6);
  assign w547[28] = |(datain[199:196] ^ 4);
  assign w547[29] = |(datain[195:192] ^ 7);
  assign w547[30] = |(datain[191:188] ^ 7);
  assign w547[31] = |(datain[187:184] ^ 5);
  assign w547[32] = |(datain[183:180] ^ 15);
  assign w547[33] = |(datain[179:176] ^ 6);
  assign comp[547] = ~(|w547);
  wire [64-1:0] w548;
  assign w548[0] = |(datain[311:308] ^ 15);
  assign w548[1] = |(datain[307:304] ^ 10);
  assign w548[2] = |(datain[303:300] ^ 12);
  assign w548[3] = |(datain[299:296] ^ 3);
  assign w548[4] = |(datain[295:292] ^ 15);
  assign w548[5] = |(datain[291:288] ^ 14);
  assign w548[6] = |(datain[287:284] ^ 8);
  assign w548[7] = |(datain[283:280] ^ 4);
  assign w548[8] = |(datain[279:276] ^ 13);
  assign w548[9] = |(datain[275:272] ^ 12);
  assign w548[10] = |(datain[271:268] ^ 0);
  assign w548[11] = |(datain[267:264] ^ 1);
  assign w548[12] = |(datain[263:260] ^ 14);
  assign w548[13] = |(datain[259:256] ^ 8);
  assign w548[14] = |(datain[255:252] ^ 14);
  assign w548[15] = |(datain[251:248] ^ 3);
  assign w548[16] = |(datain[247:244] ^ 15);
  assign w548[17] = |(datain[243:240] ^ 15);
  assign w548[18] = |(datain[239:236] ^ 11);
  assign w548[19] = |(datain[235:232] ^ 4);
  assign w548[20] = |(datain[231:228] ^ 4);
  assign w548[21] = |(datain[227:224] ^ 0);
  assign w548[22] = |(datain[223:220] ^ 8);
  assign w548[23] = |(datain[219:216] ^ 13);
  assign w548[24] = |(datain[215:212] ^ 9);
  assign w548[25] = |(datain[211:208] ^ 4);
  assign w548[26] = |(datain[207:204] ^ 0);
  assign w548[27] = |(datain[203:200] ^ 9);
  assign w548[28] = |(datain[199:196] ^ 0);
  assign w548[29] = |(datain[195:192] ^ 1);
  assign w548[30] = |(datain[191:188] ^ 11);
  assign w548[31] = |(datain[187:184] ^ 9);
  assign w548[32] = |(datain[183:180] ^ 15);
  assign w548[33] = |(datain[179:176] ^ 10);
  assign w548[34] = |(datain[175:172] ^ 0);
  assign w548[35] = |(datain[171:168] ^ 0);
  assign w548[36] = |(datain[167:164] ^ 14);
  assign w548[37] = |(datain[163:160] ^ 8);
  assign w548[38] = |(datain[159:156] ^ 0);
  assign w548[39] = |(datain[155:152] ^ 4);
  assign w548[40] = |(datain[151:148] ^ 0);
  assign w548[41] = |(datain[147:144] ^ 0);
  assign w548[42] = |(datain[143:140] ^ 14);
  assign w548[43] = |(datain[139:136] ^ 11);
  assign w548[44] = |(datain[135:132] ^ 13);
  assign w548[45] = |(datain[131:128] ^ 5);
  assign w548[46] = |(datain[127:124] ^ 11);
  assign w548[47] = |(datain[123:120] ^ 4);
  assign w548[48] = |(datain[119:116] ^ 3);
  assign w548[49] = |(datain[115:112] ^ 15);
  assign w548[50] = |(datain[111:108] ^ 8);
  assign w548[51] = |(datain[107:104] ^ 11);
  assign w548[52] = |(datain[103:100] ^ 9);
  assign w548[53] = |(datain[99:96] ^ 12);
  assign w548[54] = |(datain[95:92] ^ 0);
  assign w548[55] = |(datain[91:88] ^ 3);
  assign w548[56] = |(datain[87:84] ^ 0);
  assign w548[57] = |(datain[83:80] ^ 2);
  assign w548[58] = |(datain[79:76] ^ 12);
  assign w548[59] = |(datain[75:72] ^ 13);
  assign w548[60] = |(datain[71:68] ^ 2);
  assign w548[61] = |(datain[67:64] ^ 1);
  assign w548[62] = |(datain[63:60] ^ 12);
  assign w548[63] = |(datain[59:56] ^ 3);
  assign comp[548] = ~(|w548);
  wire [34-1:0] w549;
  assign w549[0] = |(datain[311:308] ^ 11);
  assign w549[1] = |(datain[307:304] ^ 14);
  assign w549[2] = |(datain[303:300] ^ 1);
  assign w549[3] = |(datain[299:296] ^ 6);
  assign w549[4] = |(datain[295:292] ^ 0);
  assign w549[5] = |(datain[291:288] ^ 1);
  assign w549[6] = |(datain[287:284] ^ 11);
  assign w549[7] = |(datain[283:280] ^ 9);
  assign w549[8] = |(datain[279:276] ^ 11);
  assign w549[9] = |(datain[275:272] ^ 12);
  assign w549[10] = |(datain[271:268] ^ 0);
  assign w549[11] = |(datain[267:264] ^ 1);
  assign w549[12] = |(datain[263:260] ^ 2);
  assign w549[13] = |(datain[259:256] ^ 14);
  assign w549[14] = |(datain[255:252] ^ 8);
  assign w549[15] = |(datain[251:248] ^ 1);
  assign w549[16] = |(datain[247:244] ^ 2);
  assign w549[17] = |(datain[243:240] ^ 12);
  assign w549[18] = |(datain[239:236] ^ 0);
  assign w549[19] = |(datain[235:232] ^ 0);
  assign w549[20] = |(datain[231:228] ^ 0);
  assign w549[21] = |(datain[227:224] ^ 0);
  assign w549[22] = |(datain[223:220] ^ 8);
  assign w549[23] = |(datain[219:216] ^ 3);
  assign w549[24] = |(datain[215:212] ^ 12);
  assign w549[25] = |(datain[211:208] ^ 6);
  assign w549[26] = |(datain[207:204] ^ 0);
  assign w549[27] = |(datain[203:200] ^ 2);
  assign w549[28] = |(datain[199:196] ^ 4);
  assign w549[29] = |(datain[195:192] ^ 9);
  assign w549[30] = |(datain[191:188] ^ 7);
  assign w549[31] = |(datain[187:184] ^ 5);
  assign w549[32] = |(datain[183:180] ^ 15);
  assign w549[33] = |(datain[179:176] ^ 5);
  assign comp[549] = ~(|w549);
  wire [30-1:0] w550;
  assign w550[0] = |(datain[311:308] ^ 0);
  assign w550[1] = |(datain[307:304] ^ 1);
  assign w550[2] = |(datain[303:300] ^ 11);
  assign w550[3] = |(datain[299:296] ^ 9);
  assign w550[4] = |(datain[295:292] ^ 11);
  assign w550[5] = |(datain[291:288] ^ 13);
  assign w550[6] = |(datain[287:284] ^ 0);
  assign w550[7] = |(datain[283:280] ^ 1);
  assign w550[8] = |(datain[279:276] ^ 2);
  assign w550[9] = |(datain[275:272] ^ 14);
  assign w550[10] = |(datain[271:268] ^ 8);
  assign w550[11] = |(datain[267:264] ^ 1);
  assign w550[12] = |(datain[263:260] ^ 2);
  assign w550[13] = |(datain[259:256] ^ 12);
  assign w550[14] = |(datain[255:252] ^ 0);
  assign w550[15] = |(datain[251:248] ^ 0);
  assign w550[16] = |(datain[247:244] ^ 0);
  assign w550[17] = |(datain[243:240] ^ 0);
  assign w550[18] = |(datain[239:236] ^ 8);
  assign w550[19] = |(datain[235:232] ^ 3);
  assign w550[20] = |(datain[231:228] ^ 12);
  assign w550[21] = |(datain[227:224] ^ 6);
  assign w550[22] = |(datain[223:220] ^ 0);
  assign w550[23] = |(datain[219:216] ^ 2);
  assign w550[24] = |(datain[215:212] ^ 4);
  assign w550[25] = |(datain[211:208] ^ 9);
  assign w550[26] = |(datain[207:204] ^ 7);
  assign w550[27] = |(datain[203:200] ^ 5);
  assign w550[28] = |(datain[199:196] ^ 15);
  assign w550[29] = |(datain[195:192] ^ 5);
  assign comp[550] = ~(|w550);
  wire [34-1:0] w551;
  assign w551[0] = |(datain[311:308] ^ 11);
  assign w551[1] = |(datain[307:304] ^ 11);
  assign w551[2] = |(datain[303:300] ^ 1);
  assign w551[3] = |(datain[299:296] ^ 4);
  assign w551[4] = |(datain[295:292] ^ 0);
  assign w551[5] = |(datain[291:288] ^ 1);
  assign w551[6] = |(datain[287:284] ^ 11);
  assign w551[7] = |(datain[283:280] ^ 9);
  assign w551[8] = |(datain[279:276] ^ 13);
  assign w551[9] = |(datain[275:272] ^ 10);
  assign w551[10] = |(datain[271:268] ^ 0);
  assign w551[11] = |(datain[267:264] ^ 1);
  assign w551[12] = |(datain[263:260] ^ 2);
  assign w551[13] = |(datain[259:256] ^ 14);
  assign w551[14] = |(datain[255:252] ^ 8);
  assign w551[15] = |(datain[251:248] ^ 1);
  assign w551[16] = |(datain[247:244] ^ 3);
  assign w551[17] = |(datain[243:240] ^ 7);
  assign w551[18] = |(datain[239:236] ^ 0);
  assign w551[19] = |(datain[235:232] ^ 0);
  assign w551[20] = |(datain[231:228] ^ 0);
  assign w551[21] = |(datain[227:224] ^ 0);
  assign w551[22] = |(datain[223:220] ^ 8);
  assign w551[23] = |(datain[219:216] ^ 3);
  assign w551[24] = |(datain[215:212] ^ 12);
  assign w551[25] = |(datain[211:208] ^ 3);
  assign w551[26] = |(datain[207:204] ^ 0);
  assign w551[27] = |(datain[203:200] ^ 2);
  assign w551[28] = |(datain[199:196] ^ 4);
  assign w551[29] = |(datain[195:192] ^ 9);
  assign w551[30] = |(datain[191:188] ^ 7);
  assign w551[31] = |(datain[187:184] ^ 5);
  assign w551[32] = |(datain[183:180] ^ 15);
  assign w551[33] = |(datain[179:176] ^ 5);
  assign comp[551] = ~(|w551);
  wire [42-1:0] w552;
  assign w552[0] = |(datain[311:308] ^ 0);
  assign w552[1] = |(datain[307:304] ^ 5);
  assign w552[2] = |(datain[303:300] ^ 0);
  assign w552[3] = |(datain[299:296] ^ 0);
  assign w552[4] = |(datain[295:292] ^ 8);
  assign w552[5] = |(datain[291:288] ^ 10);
  assign w552[6] = |(datain[287:284] ^ 2);
  assign w552[7] = |(datain[283:280] ^ 5);
  assign w552[8] = |(datain[279:276] ^ 3);
  assign w552[9] = |(datain[275:272] ^ 10);
  assign w552[10] = |(datain[271:268] ^ 2);
  assign w552[11] = |(datain[267:264] ^ 4);
  assign w552[12] = |(datain[263:260] ^ 7);
  assign w552[13] = |(datain[259:256] ^ 5);
  assign w552[14] = |(datain[255:252] ^ 0);
  assign w552[15] = |(datain[251:248] ^ 7);
  assign w552[16] = |(datain[247:244] ^ 4);
  assign w552[17] = |(datain[243:240] ^ 6);
  assign w552[18] = |(datain[239:236] ^ 4);
  assign w552[19] = |(datain[235:232] ^ 7);
  assign w552[20] = |(datain[231:228] ^ 14);
  assign w552[21] = |(datain[227:224] ^ 2);
  assign w552[22] = |(datain[223:220] ^ 15);
  assign w552[23] = |(datain[219:216] ^ 6);
  assign w552[24] = |(datain[215:212] ^ 14);
  assign w552[25] = |(datain[211:208] ^ 11);
  assign w552[26] = |(datain[207:204] ^ 7);
  assign w552[27] = |(datain[203:200] ^ 2);
  assign w552[28] = |(datain[199:196] ^ 9);
  assign w552[29] = |(datain[195:192] ^ 0);
  assign w552[30] = |(datain[191:188] ^ 5);
  assign w552[31] = |(datain[187:184] ^ 14);
  assign w552[32] = |(datain[183:180] ^ 11);
  assign w552[33] = |(datain[179:176] ^ 8);
  assign w552[34] = |(datain[175:172] ^ 0);
  assign w552[35] = |(datain[171:168] ^ 0);
  assign w552[36] = |(datain[167:164] ^ 4);
  assign w552[37] = |(datain[163:160] ^ 2);
  assign w552[38] = |(datain[159:156] ^ 8);
  assign w552[39] = |(datain[155:152] ^ 11);
  assign w552[40] = |(datain[151:148] ^ 9);
  assign w552[41] = |(datain[147:144] ^ 12);
  assign comp[552] = ~(|w552);
  wire [44-1:0] w553;
  assign w553[0] = |(datain[311:308] ^ 9);
  assign w553[1] = |(datain[307:304] ^ 9);
  assign w553[2] = |(datain[303:300] ^ 7);
  assign w553[3] = |(datain[299:296] ^ 5);
  assign w553[4] = |(datain[295:292] ^ 0);
  assign w553[5] = |(datain[291:288] ^ 2);
  assign w553[6] = |(datain[287:284] ^ 9);
  assign w553[7] = |(datain[283:280] ^ 3);
  assign w553[8] = |(datain[279:276] ^ 12);
  assign w553[9] = |(datain[275:272] ^ 15);
  assign w553[10] = |(datain[271:268] ^ 9);
  assign w553[11] = |(datain[267:264] ^ 12);
  assign w553[12] = |(datain[263:260] ^ 3);
  assign w553[13] = |(datain[259:256] ^ 13);
  assign w553[14] = |(datain[255:252] ^ 0);
  assign w553[15] = |(datain[251:248] ^ 0);
  assign w553[16] = |(datain[247:244] ^ 4);
  assign w553[17] = |(datain[243:240] ^ 11);
  assign w553[18] = |(datain[239:236] ^ 7);
  assign w553[19] = |(datain[235:232] ^ 5);
  assign w553[20] = |(datain[231:228] ^ 6);
  assign w553[21] = |(datain[227:224] ^ 1);
  assign w553[22] = |(datain[223:220] ^ 6);
  assign w553[23] = |(datain[219:216] ^ 0);
  assign w553[24] = |(datain[215:212] ^ 1);
  assign w553[25] = |(datain[211:208] ^ 14);
  assign w553[26] = |(datain[207:204] ^ 0);
  assign w553[27] = |(datain[203:200] ^ 6);
  assign w553[28] = |(datain[199:196] ^ 11);
  assign w553[29] = |(datain[195:192] ^ 0);
  assign w553[30] = |(datain[191:188] ^ 0);
  assign w553[31] = |(datain[187:184] ^ 1);
  assign w553[32] = |(datain[183:180] ^ 3);
  assign w553[33] = |(datain[179:176] ^ 3);
  assign w553[34] = |(datain[175:172] ^ 12);
  assign w553[35] = |(datain[171:168] ^ 9);
  assign w553[36] = |(datain[167:164] ^ 11);
  assign w553[37] = |(datain[163:160] ^ 4);
  assign w553[38] = |(datain[159:156] ^ 4);
  assign w553[39] = |(datain[155:152] ^ 3);
  assign w553[40] = |(datain[151:148] ^ 12);
  assign w553[41] = |(datain[147:144] ^ 13);
  assign w553[42] = |(datain[143:140] ^ 2);
  assign w553[43] = |(datain[139:136] ^ 1);
  assign comp[553] = ~(|w553);
  wire [76-1:0] w554;
  assign w554[0] = |(datain[311:308] ^ 0);
  assign w554[1] = |(datain[307:304] ^ 6);
  assign w554[2] = |(datain[303:300] ^ 11);
  assign w554[3] = |(datain[299:296] ^ 6);
  assign w554[4] = |(datain[295:292] ^ 0);
  assign w554[5] = |(datain[291:288] ^ 5);
  assign w554[6] = |(datain[287:284] ^ 14);
  assign w554[7] = |(datain[283:280] ^ 9);
  assign w554[8] = |(datain[279:276] ^ 2);
  assign w554[9] = |(datain[275:272] ^ 14);
  assign w554[10] = |(datain[271:268] ^ 10);
  assign w554[11] = |(datain[267:264] ^ 1);
  assign w554[12] = |(datain[263:260] ^ 2);
  assign w554[13] = |(datain[259:256] ^ 0);
  assign w554[14] = |(datain[255:252] ^ 0);
  assign w554[15] = |(datain[251:248] ^ 1);
  assign w554[16] = |(datain[247:244] ^ 2);
  assign w554[17] = |(datain[243:240] ^ 13);
  assign w554[18] = |(datain[239:236] ^ 0);
  assign w554[19] = |(datain[235:232] ^ 3);
  assign w554[20] = |(datain[231:228] ^ 0);
  assign w554[21] = |(datain[227:224] ^ 0);
  assign w554[22] = |(datain[223:220] ^ 10);
  assign w554[23] = |(datain[219:216] ^ 3);
  assign w554[24] = |(datain[215:212] ^ 11);
  assign w554[25] = |(datain[211:208] ^ 7);
  assign w554[26] = |(datain[207:204] ^ 0);
  assign w554[27] = |(datain[203:200] ^ 5);
  assign w554[28] = |(datain[199:196] ^ 11);
  assign w554[29] = |(datain[195:192] ^ 8);
  assign w554[30] = |(datain[191:188] ^ 0);
  assign w554[31] = |(datain[187:184] ^ 0);
  assign w554[32] = |(datain[183:180] ^ 4);
  assign w554[33] = |(datain[179:176] ^ 2);
  assign w554[34] = |(datain[175:172] ^ 3);
  assign w554[35] = |(datain[171:168] ^ 3);
  assign w554[36] = |(datain[167:164] ^ 12);
  assign w554[37] = |(datain[163:160] ^ 9);
  assign w554[38] = |(datain[159:156] ^ 3);
  assign w554[39] = |(datain[155:152] ^ 3);
  assign w554[40] = |(datain[151:148] ^ 13);
  assign w554[41] = |(datain[147:144] ^ 2);
  assign w554[42] = |(datain[143:140] ^ 12);
  assign w554[43] = |(datain[139:136] ^ 13);
  assign w554[44] = |(datain[135:132] ^ 2);
  assign w554[45] = |(datain[131:128] ^ 1);
  assign w554[46] = |(datain[127:124] ^ 7);
  assign w554[47] = |(datain[123:120] ^ 2);
  assign w554[48] = |(datain[119:116] ^ 0);
  assign w554[49] = |(datain[115:112] ^ 10);
  assign w554[50] = |(datain[111:108] ^ 11);
  assign w554[51] = |(datain[107:104] ^ 4);
  assign w554[52] = |(datain[103:100] ^ 4);
  assign w554[53] = |(datain[99:96] ^ 0);
  assign w554[54] = |(datain[95:92] ^ 11);
  assign w554[55] = |(datain[91:88] ^ 9);
  assign w554[56] = |(datain[87:84] ^ 0);
  assign w554[57] = |(datain[83:80] ^ 3);
  assign w554[58] = |(datain[79:76] ^ 0);
  assign w554[59] = |(datain[75:72] ^ 0);
  assign w554[60] = |(datain[71:68] ^ 11);
  assign w554[61] = |(datain[67:64] ^ 10);
  assign w554[62] = |(datain[63:60] ^ 11);
  assign w554[63] = |(datain[59:56] ^ 6);
  assign w554[64] = |(datain[55:52] ^ 0);
  assign w554[65] = |(datain[51:48] ^ 5);
  assign w554[66] = |(datain[47:44] ^ 12);
  assign w554[67] = |(datain[43:40] ^ 13);
  assign w554[68] = |(datain[39:36] ^ 2);
  assign w554[69] = |(datain[35:32] ^ 1);
  assign w554[70] = |(datain[31:28] ^ 11);
  assign w554[71] = |(datain[27:24] ^ 8);
  assign w554[72] = |(datain[23:20] ^ 0);
  assign w554[73] = |(datain[19:16] ^ 1);
  assign w554[74] = |(datain[15:12] ^ 5);
  assign w554[75] = |(datain[11:8] ^ 7);
  assign comp[554] = ~(|w554);
  wire [30-1:0] w555;
  assign w555[0] = |(datain[311:308] ^ 1);
  assign w555[1] = |(datain[307:304] ^ 14);
  assign w555[2] = |(datain[303:300] ^ 7);
  assign w555[3] = |(datain[299:296] ^ 1);
  assign w555[4] = |(datain[295:292] ^ 0);
  assign w555[5] = |(datain[291:288] ^ 5);
  assign w555[6] = |(datain[287:284] ^ 11);
  assign w555[7] = |(datain[283:280] ^ 10);
  assign w555[8] = |(datain[279:276] ^ 14);
  assign w555[9] = |(datain[275:272] ^ 1);
  assign w555[10] = |(datain[271:268] ^ 0);
  assign w555[11] = |(datain[267:264] ^ 3);
  assign w555[12] = |(datain[263:260] ^ 11);
  assign w555[13] = |(datain[259:256] ^ 8);
  assign w555[14] = |(datain[255:252] ^ 0);
  assign w555[15] = |(datain[251:248] ^ 0);
  assign w555[16] = |(datain[247:244] ^ 3);
  assign w555[17] = |(datain[243:240] ^ 13);
  assign w555[18] = |(datain[239:236] ^ 12);
  assign w555[19] = |(datain[235:232] ^ 13);
  assign w555[20] = |(datain[231:228] ^ 2);
  assign w555[21] = |(datain[227:224] ^ 1);
  assign w555[22] = |(datain[223:220] ^ 7);
  assign w555[23] = |(datain[219:216] ^ 2);
  assign w555[24] = |(datain[215:212] ^ 3);
  assign w555[25] = |(datain[211:208] ^ 3);
  assign w555[26] = |(datain[207:204] ^ 8);
  assign w555[27] = |(datain[203:200] ^ 11);
  assign w555[28] = |(datain[199:196] ^ 13);
  assign w555[29] = |(datain[195:192] ^ 8);
  assign comp[555] = ~(|w555);
  wire [44-1:0] w556;
  assign w556[0] = |(datain[311:308] ^ 11);
  assign w556[1] = |(datain[307:304] ^ 4);
  assign w556[2] = |(datain[303:300] ^ 2);
  assign w556[3] = |(datain[299:296] ^ 10);
  assign w556[4] = |(datain[295:292] ^ 12);
  assign w556[5] = |(datain[291:288] ^ 13);
  assign w556[6] = |(datain[287:284] ^ 2);
  assign w556[7] = |(datain[283:280] ^ 1);
  assign w556[8] = |(datain[279:276] ^ 8);
  assign w556[9] = |(datain[275:272] ^ 1);
  assign w556[10] = |(datain[271:268] ^ 15);
  assign w556[11] = |(datain[267:264] ^ 10);
  assign w556[12] = |(datain[263:260] ^ 1);
  assign w556[13] = |(datain[259:256] ^ 9);
  assign w556[14] = |(datain[255:252] ^ 0);
  assign w556[15] = |(datain[251:248] ^ 5);
  assign w556[16] = |(datain[247:244] ^ 7);
  assign w556[17] = |(datain[243:240] ^ 4);
  assign w556[18] = |(datain[239:236] ^ 1);
  assign w556[19] = |(datain[235:232] ^ 5);
  assign w556[20] = |(datain[231:228] ^ 8);
  assign w556[21] = |(datain[227:224] ^ 1);
  assign w556[22] = |(datain[223:220] ^ 15);
  assign w556[23] = |(datain[219:216] ^ 10);
  assign w556[24] = |(datain[215:212] ^ 1);
  assign w556[25] = |(datain[211:208] ^ 4);
  assign w556[26] = |(datain[207:204] ^ 0);
  assign w556[27] = |(datain[203:200] ^ 6);
  assign w556[28] = |(datain[199:196] ^ 7);
  assign w556[29] = |(datain[195:192] ^ 4);
  assign w556[30] = |(datain[191:188] ^ 1);
  assign w556[31] = |(datain[187:184] ^ 5);
  assign w556[32] = |(datain[183:180] ^ 8);
  assign w556[33] = |(datain[179:176] ^ 1);
  assign w556[34] = |(datain[175:172] ^ 15);
  assign w556[35] = |(datain[171:168] ^ 10);
  assign w556[36] = |(datain[167:164] ^ 0);
  assign w556[37] = |(datain[163:160] ^ 9);
  assign w556[38] = |(datain[159:156] ^ 0);
  assign w556[39] = |(datain[155:152] ^ 7);
  assign w556[40] = |(datain[151:148] ^ 7);
  assign w556[41] = |(datain[147:144] ^ 4);
  assign w556[42] = |(datain[143:140] ^ 1);
  assign w556[43] = |(datain[139:136] ^ 5);
  assign comp[556] = ~(|w556);
  wire [32-1:0] w557;
  assign w557[0] = |(datain[311:308] ^ 8);
  assign w557[1] = |(datain[307:304] ^ 1);
  assign w557[2] = |(datain[303:300] ^ 14);
  assign w557[3] = |(datain[299:296] ^ 9);
  assign w557[4] = |(datain[295:292] ^ 14);
  assign w557[5] = |(datain[291:288] ^ 1);
  assign w557[6] = |(datain[287:284] ^ 0);
  assign w557[7] = |(datain[283:280] ^ 5);
  assign w557[8] = |(datain[279:276] ^ 11);
  assign w557[9] = |(datain[275:272] ^ 4);
  assign w557[10] = |(datain[271:268] ^ 15);
  assign w557[11] = |(datain[267:264] ^ 10);
  assign w557[12] = |(datain[263:260] ^ 12);
  assign w557[13] = |(datain[259:256] ^ 13);
  assign w557[14] = |(datain[255:252] ^ 2);
  assign w557[15] = |(datain[251:248] ^ 1);
  assign w557[16] = |(datain[247:244] ^ 11);
  assign w557[17] = |(datain[243:240] ^ 8);
  assign w557[18] = |(datain[239:236] ^ 2);
  assign w557[19] = |(datain[235:232] ^ 1);
  assign w557[20] = |(datain[231:228] ^ 3);
  assign w557[21] = |(datain[227:224] ^ 5);
  assign w557[22] = |(datain[223:220] ^ 12);
  assign w557[23] = |(datain[219:216] ^ 13);
  assign w557[24] = |(datain[215:212] ^ 2);
  assign w557[25] = |(datain[211:208] ^ 1);
  assign w557[26] = |(datain[207:204] ^ 8);
  assign w557[27] = |(datain[203:200] ^ 9);
  assign w557[28] = |(datain[199:196] ^ 1);
  assign w557[29] = |(datain[195:192] ^ 14);
  assign w557[30] = |(datain[191:188] ^ 1);
  assign w557[31] = |(datain[187:184] ^ 10);
  assign comp[557] = ~(|w557);
  wire [42-1:0] w558;
  assign w558[0] = |(datain[311:308] ^ 5);
  assign w558[1] = |(datain[307:304] ^ 14);
  assign w558[2] = |(datain[303:300] ^ 1);
  assign w558[3] = |(datain[299:296] ^ 14);
  assign w558[4] = |(datain[295:292] ^ 0);
  assign w558[5] = |(datain[291:288] ^ 14);
  assign w558[6] = |(datain[287:284] ^ 0);
  assign w558[7] = |(datain[283:280] ^ 14);
  assign w558[8] = |(datain[279:276] ^ 0);
  assign w558[9] = |(datain[275:272] ^ 7);
  assign w558[10] = |(datain[271:268] ^ 1);
  assign w558[11] = |(datain[267:264] ^ 15);
  assign w558[12] = |(datain[263:260] ^ 11);
  assign w558[13] = |(datain[259:256] ^ 9);
  assign w558[14] = |(datain[255:252] ^ 15);
  assign w558[15] = |(datain[251:248] ^ 6);
  assign w558[16] = |(datain[247:244] ^ 0);
  assign w558[17] = |(datain[243:240] ^ 10);
  assign w558[18] = |(datain[239:236] ^ 8);
  assign w558[19] = |(datain[235:232] ^ 3);
  assign w558[20] = |(datain[231:228] ^ 14);
  assign w558[21] = |(datain[227:224] ^ 14);
  assign w558[22] = |(datain[223:220] ^ 0);
  assign w558[23] = |(datain[219:216] ^ 4);
  assign w558[24] = |(datain[215:212] ^ 8);
  assign w558[25] = |(datain[211:208] ^ 11);
  assign w558[26] = |(datain[207:204] ^ 15);
  assign w558[27] = |(datain[203:200] ^ 14);
  assign w558[28] = |(datain[199:196] ^ 15);
  assign w558[29] = |(datain[195:192] ^ 13);
  assign w558[30] = |(datain[191:188] ^ 10);
  assign w558[31] = |(datain[187:184] ^ 12);
  assign w558[32] = |(datain[183:180] ^ 3);
  assign w558[33] = |(datain[179:176] ^ 4);
  assign w558[34] = |(datain[175:172] ^ 15);
  assign w558[35] = |(datain[171:168] ^ 6);
  assign w558[36] = |(datain[167:164] ^ 10);
  assign w558[37] = |(datain[163:160] ^ 10);
  assign w558[38] = |(datain[159:156] ^ 14);
  assign w558[39] = |(datain[155:152] ^ 2);
  assign w558[40] = |(datain[151:148] ^ 15);
  assign w558[41] = |(datain[147:144] ^ 10);
  assign comp[558] = ~(|w558);
  wire [42-1:0] w559;
  assign w559[0] = |(datain[311:308] ^ 15);
  assign w559[1] = |(datain[307:304] ^ 12);
  assign w559[2] = |(datain[303:300] ^ 3);
  assign w559[3] = |(datain[299:296] ^ 6);
  assign w559[4] = |(datain[295:292] ^ 8);
  assign w559[5] = |(datain[291:288] ^ 10);
  assign w559[6] = |(datain[287:284] ^ 4);
  assign w559[7] = |(datain[283:280] ^ 5);
  assign w559[8] = |(datain[279:276] ^ 13);
  assign w559[9] = |(datain[275:272] ^ 4);
  assign w559[10] = |(datain[271:268] ^ 2);
  assign w559[11] = |(datain[267:264] ^ 8);
  assign w559[12] = |(datain[263:260] ^ 4);
  assign w559[13] = |(datain[259:256] ^ 6);
  assign w559[14] = |(datain[255:252] ^ 0);
  assign w559[15] = |(datain[251:248] ^ 0);
  assign w559[16] = |(datain[247:244] ^ 8);
  assign w559[17] = |(datain[243:240] ^ 0);
  assign w559[18] = |(datain[239:236] ^ 4);
  assign w559[19] = |(datain[235:232] ^ 6);
  assign w559[20] = |(datain[231:228] ^ 0);
  assign w559[21] = |(datain[227:224] ^ 0);
  assign w559[22] = |(datain[223:220] ^ 15);
  assign w559[23] = |(datain[219:216] ^ 2);
  assign w559[24] = |(datain[215:212] ^ 4);
  assign w559[25] = |(datain[211:208] ^ 9);
  assign w559[26] = |(datain[207:204] ^ 7);
  assign w559[27] = |(datain[203:200] ^ 8);
  assign w559[28] = |(datain[199:196] ^ 0);
  assign w559[29] = |(datain[195:192] ^ 6);
  assign w559[30] = |(datain[191:188] ^ 4);
  assign w559[31] = |(datain[187:184] ^ 13);
  assign w559[32] = |(datain[183:180] ^ 4);
  assign w559[33] = |(datain[179:176] ^ 14);
  assign w559[34] = |(datain[175:172] ^ 7);
  assign w559[35] = |(datain[171:168] ^ 9);
  assign w559[36] = |(datain[167:164] ^ 14);
  assign w559[37] = |(datain[163:160] ^ 10);
  assign w559[38] = |(datain[159:156] ^ 14);
  assign w559[39] = |(datain[155:152] ^ 11);
  assign w559[40] = |(datain[151:148] ^ 14);
  assign w559[41] = |(datain[147:144] ^ 5);
  assign comp[559] = ~(|w559);
  wire [44-1:0] w560;
  assign w560[0] = |(datain[311:308] ^ 14);
  assign w560[1] = |(datain[307:304] ^ 12);
  assign w560[2] = |(datain[303:300] ^ 8);
  assign w560[3] = |(datain[299:296] ^ 3);
  assign w560[4] = |(datain[295:292] ^ 12);
  assign w560[5] = |(datain[291:288] ^ 4);
  assign w560[6] = |(datain[287:284] ^ 14);
  assign w560[7] = |(datain[283:280] ^ 14);
  assign w560[8] = |(datain[279:276] ^ 14);
  assign w560[9] = |(datain[275:272] ^ 8);
  assign w560[10] = |(datain[271:268] ^ 8);
  assign w560[11] = |(datain[267:264] ^ 3);
  assign w560[12] = |(datain[263:260] ^ 0);
  assign w560[13] = |(datain[259:256] ^ 3);
  assign w560[14] = |(datain[255:252] ^ 11);
  assign w560[15] = |(datain[251:248] ^ 8);
  assign w560[16] = |(datain[247:244] ^ 11);
  assign w560[17] = |(datain[243:240] ^ 6);
  assign w560[18] = |(datain[239:236] ^ 1);
  assign w560[19] = |(datain[235:232] ^ 4);
  assign w560[20] = |(datain[231:228] ^ 5);
  assign w560[21] = |(datain[227:224] ^ 0);
  assign w560[22] = |(datain[223:220] ^ 14);
  assign w560[23] = |(datain[219:216] ^ 8);
  assign w560[24] = |(datain[215:212] ^ 3);
  assign w560[25] = |(datain[211:208] ^ 14);
  assign w560[26] = |(datain[207:204] ^ 0);
  assign w560[27] = |(datain[203:200] ^ 11);
  assign w560[28] = |(datain[199:196] ^ 5);
  assign w560[29] = |(datain[195:192] ^ 0);
  assign w560[30] = |(datain[191:188] ^ 14);
  assign w560[31] = |(datain[187:184] ^ 8);
  assign w560[32] = |(datain[183:180] ^ 4);
  assign w560[33] = |(datain[179:176] ^ 5);
  assign w560[34] = |(datain[175:172] ^ 0);
  assign w560[35] = |(datain[171:168] ^ 11);
  assign w560[36] = |(datain[167:164] ^ 8);
  assign w560[37] = |(datain[163:160] ^ 3);
  assign w560[38] = |(datain[159:156] ^ 12);
  assign w560[39] = |(datain[155:152] ^ 4);
  assign w560[40] = |(datain[151:148] ^ 0);
  assign w560[41] = |(datain[147:144] ^ 4);
  assign w560[42] = |(datain[143:140] ^ 11);
  assign w560[43] = |(datain[139:136] ^ 8);
  assign comp[560] = ~(|w560);
  wire [76-1:0] w561;
  assign w561[0] = |(datain[311:308] ^ 11);
  assign w561[1] = |(datain[307:304] ^ 9);
  assign w561[2] = |(datain[303:300] ^ 3);
  assign w561[3] = |(datain[299:296] ^ 11);
  assign w561[4] = |(datain[295:292] ^ 0);
  assign w561[5] = |(datain[291:288] ^ 0);
  assign w561[6] = |(datain[287:284] ^ 8);
  assign w561[7] = |(datain[283:280] ^ 13);
  assign w561[8] = |(datain[279:276] ^ 9);
  assign w561[9] = |(datain[275:272] ^ 4);
  assign w561[10] = |(datain[271:268] ^ 15);
  assign w561[11] = |(datain[267:264] ^ 4);
  assign w561[12] = |(datain[263:260] ^ 0);
  assign w561[13] = |(datain[259:256] ^ 0);
  assign w561[14] = |(datain[255:252] ^ 12);
  assign w561[15] = |(datain[251:248] ^ 13);
  assign w561[16] = |(datain[247:244] ^ 2);
  assign w561[17] = |(datain[243:240] ^ 1);
  assign w561[18] = |(datain[239:236] ^ 8);
  assign w561[19] = |(datain[235:232] ^ 13);
  assign w561[20] = |(datain[231:228] ^ 9);
  assign w561[21] = |(datain[227:224] ^ 4);
  assign w561[22] = |(datain[223:220] ^ 2);
  assign w561[23] = |(datain[219:216] ^ 0);
  assign w561[24] = |(datain[215:212] ^ 0);
  assign w561[25] = |(datain[211:208] ^ 2);
  assign w561[26] = |(datain[207:204] ^ 11);
  assign w561[27] = |(datain[203:200] ^ 9);
  assign w561[28] = |(datain[199:196] ^ 15);
  assign w561[29] = |(datain[195:192] ^ 1);
  assign w561[30] = |(datain[191:188] ^ 0);
  assign w561[31] = |(datain[187:184] ^ 1);
  assign w561[32] = |(datain[183:180] ^ 11);
  assign w561[33] = |(datain[179:176] ^ 4);
  assign w561[34] = |(datain[175:172] ^ 4);
  assign w561[35] = |(datain[171:168] ^ 0);
  assign w561[36] = |(datain[167:164] ^ 12);
  assign w561[37] = |(datain[163:160] ^ 13);
  assign w561[38] = |(datain[159:156] ^ 2);
  assign w561[39] = |(datain[155:152] ^ 1);
  assign w561[40] = |(datain[151:148] ^ 14);
  assign w561[41] = |(datain[147:144] ^ 4);
  assign w561[42] = |(datain[143:140] ^ 4);
  assign w561[43] = |(datain[139:136] ^ 0);
  assign w561[44] = |(datain[135:132] ^ 8);
  assign w561[45] = |(datain[131:128] ^ 10);
  assign w561[46] = |(datain[127:124] ^ 12);
  assign w561[47] = |(datain[123:120] ^ 8);
  assign w561[48] = |(datain[119:116] ^ 3);
  assign w561[49] = |(datain[115:112] ^ 2);
  assign w561[50] = |(datain[111:108] ^ 14);
  assign w561[51] = |(datain[107:104] ^ 13);
  assign w561[52] = |(datain[103:100] ^ 14);
  assign w561[53] = |(datain[99:96] ^ 4);
  assign w561[54] = |(datain[95:92] ^ 4);
  assign w561[55] = |(datain[91:88] ^ 0);
  assign w561[56] = |(datain[87:84] ^ 3);
  assign w561[57] = |(datain[83:80] ^ 2);
  assign w561[58] = |(datain[79:76] ^ 12);
  assign w561[59] = |(datain[75:72] ^ 8);
  assign w561[60] = |(datain[71:68] ^ 14);
  assign w561[61] = |(datain[67:64] ^ 5);
  assign w561[62] = |(datain[63:60] ^ 4);
  assign w561[63] = |(datain[59:56] ^ 0);
  assign w561[64] = |(datain[55:52] ^ 8);
  assign w561[65] = |(datain[51:48] ^ 11);
  assign w561[66] = |(datain[47:44] ^ 13);
  assign w561[67] = |(datain[43:40] ^ 0);
  assign w561[68] = |(datain[39:36] ^ 14);
  assign w561[69] = |(datain[35:32] ^ 5);
  assign w561[70] = |(datain[31:28] ^ 4);
  assign w561[71] = |(datain[27:24] ^ 0);
  assign w561[72] = |(datain[23:20] ^ 3);
  assign w561[73] = |(datain[19:16] ^ 3);
  assign w561[74] = |(datain[15:12] ^ 12);
  assign w561[75] = |(datain[11:8] ^ 2);
  assign comp[561] = ~(|w561);
  wire [76-1:0] w562;
  assign w562[0] = |(datain[311:308] ^ 14);
  assign w562[1] = |(datain[307:304] ^ 9);
  assign w562[2] = |(datain[303:300] ^ 3);
  assign w562[3] = |(datain[299:296] ^ 1);
  assign w562[4] = |(datain[295:292] ^ 0);
  assign w562[5] = |(datain[291:288] ^ 0);
  assign w562[6] = |(datain[287:284] ^ 5);
  assign w562[7] = |(datain[283:280] ^ 14);
  assign w562[8] = |(datain[279:276] ^ 14);
  assign w562[9] = |(datain[275:272] ^ 8);
  assign w562[10] = |(datain[271:268] ^ 0);
  assign w562[11] = |(datain[267:264] ^ 0);
  assign w562[12] = |(datain[263:260] ^ 0);
  assign w562[13] = |(datain[259:256] ^ 0);
  assign w562[14] = |(datain[255:252] ^ 5);
  assign w562[15] = |(datain[251:248] ^ 14);
  assign w562[16] = |(datain[247:244] ^ 11);
  assign w562[17] = |(datain[243:240] ^ 9);
  assign w562[18] = |(datain[239:236] ^ 15);
  assign w562[19] = |(datain[235:232] ^ 5);
  assign w562[20] = |(datain[231:228] ^ 0);
  assign w562[21] = |(datain[227:224] ^ 1);
  assign w562[22] = |(datain[223:220] ^ 8);
  assign w562[23] = |(datain[219:216] ^ 13);
  assign w562[24] = |(datain[215:212] ^ 9);
  assign w562[25] = |(datain[211:208] ^ 12);
  assign w562[26] = |(datain[207:204] ^ 2);
  assign w562[27] = |(datain[203:200] ^ 13);
  assign w562[28] = |(datain[199:196] ^ 0);
  assign w562[29] = |(datain[195:192] ^ 0);
  assign w562[30] = |(datain[191:188] ^ 11);
  assign w562[31] = |(datain[187:184] ^ 4);
  assign w562[32] = |(datain[183:180] ^ 0);
  assign w562[33] = |(datain[179:176] ^ 0);
  assign w562[34] = |(datain[175:172] ^ 2);
  assign w562[35] = |(datain[171:168] ^ 14);
  assign w562[36] = |(datain[167:164] ^ 8);
  assign w562[37] = |(datain[163:160] ^ 10);
  assign w562[38] = |(datain[159:156] ^ 0);
  assign w562[39] = |(datain[155:152] ^ 7);
  assign w562[40] = |(datain[151:148] ^ 3);
  assign w562[41] = |(datain[147:144] ^ 2);
  assign w562[42] = |(datain[143:140] ^ 12);
  assign w562[43] = |(datain[139:136] ^ 4);
  assign w562[44] = |(datain[135:132] ^ 2);
  assign w562[45] = |(datain[131:128] ^ 14);
  assign w562[46] = |(datain[127:124] ^ 8);
  assign w562[47] = |(datain[123:120] ^ 8);
  assign w562[48] = |(datain[119:116] ^ 0);
  assign w562[49] = |(datain[115:112] ^ 7);
  assign w562[50] = |(datain[111:108] ^ 14);
  assign w562[51] = |(datain[107:104] ^ 8);
  assign w562[52] = |(datain[103:100] ^ 0);
  assign w562[53] = |(datain[99:96] ^ 14);
  assign w562[54] = |(datain[95:92] ^ 0);
  assign w562[55] = |(datain[91:88] ^ 0);
  assign w562[56] = |(datain[87:84] ^ 7);
  assign w562[57] = |(datain[83:80] ^ 4);
  assign w562[58] = |(datain[79:76] ^ 0);
  assign w562[59] = |(datain[75:72] ^ 3);
  assign w562[60] = |(datain[71:68] ^ 14);
  assign w562[61] = |(datain[67:64] ^ 9);
  assign w562[62] = |(datain[63:60] ^ 1);
  assign w562[63] = |(datain[59:56] ^ 3);
  assign w562[64] = |(datain[55:52] ^ 0);
  assign w562[65] = |(datain[51:48] ^ 0);
  assign w562[66] = |(datain[47:44] ^ 4);
  assign w562[67] = |(datain[43:40] ^ 3);
  assign w562[68] = |(datain[39:36] ^ 8);
  assign w562[69] = |(datain[35:32] ^ 0);
  assign w562[70] = |(datain[31:28] ^ 12);
  assign w562[71] = |(datain[27:24] ^ 4);
  assign w562[72] = |(datain[23:20] ^ 0);
  assign w562[73] = |(datain[19:16] ^ 5);
  assign w562[74] = |(datain[15:12] ^ 14);
  assign w562[75] = |(datain[11:8] ^ 2);
  assign comp[562] = ~(|w562);
  wire [76-1:0] w563;
  assign w563[0] = |(datain[311:308] ^ 0);
  assign w563[1] = |(datain[307:304] ^ 14);
  assign w563[2] = |(datain[303:300] ^ 1);
  assign w563[3] = |(datain[299:296] ^ 7);
  assign w563[4] = |(datain[295:292] ^ 9);
  assign w563[5] = |(datain[291:288] ^ 12);
  assign w563[6] = |(datain[287:284] ^ 5);
  assign w563[7] = |(datain[283:280] ^ 8);
  assign w563[8] = |(datain[279:276] ^ 15);
  assign w563[9] = |(datain[275:272] ^ 6);
  assign w563[10] = |(datain[271:268] ^ 12);
  assign w563[11] = |(datain[267:264] ^ 4);
  assign w563[12] = |(datain[263:260] ^ 0);
  assign w563[13] = |(datain[259:256] ^ 1);
  assign w563[14] = |(datain[255:252] ^ 7);
  assign w563[15] = |(datain[251:248] ^ 4);
  assign w563[16] = |(datain[247:244] ^ 0);
  assign w563[17] = |(datain[243:240] ^ 3);
  assign w563[18] = |(datain[239:236] ^ 14);
  assign w563[19] = |(datain[235:232] ^ 11);
  assign w563[20] = |(datain[231:228] ^ 3);
  assign w563[21] = |(datain[227:224] ^ 3);
  assign w563[22] = |(datain[223:220] ^ 9);
  assign w563[23] = |(datain[219:216] ^ 0);
  assign w563[24] = |(datain[215:212] ^ 5);
  assign w563[25] = |(datain[211:208] ^ 14);
  assign w563[26] = |(datain[207:204] ^ 14);
  assign w563[27] = |(datain[203:200] ^ 8);
  assign w563[28] = |(datain[199:196] ^ 0);
  assign w563[29] = |(datain[195:192] ^ 0);
  assign w563[30] = |(datain[191:188] ^ 0);
  assign w563[31] = |(datain[187:184] ^ 0);
  assign w563[32] = |(datain[183:180] ^ 5);
  assign w563[33] = |(datain[179:176] ^ 14);
  assign w563[34] = |(datain[175:172] ^ 11);
  assign w563[35] = |(datain[171:168] ^ 9);
  assign w563[36] = |(datain[167:164] ^ 15);
  assign w563[37] = |(datain[163:160] ^ 9);
  assign w563[38] = |(datain[159:156] ^ 0);
  assign w563[39] = |(datain[155:152] ^ 1);
  assign w563[40] = |(datain[151:148] ^ 9);
  assign w563[41] = |(datain[147:144] ^ 0);
  assign w563[42] = |(datain[143:140] ^ 8);
  assign w563[43] = |(datain[139:136] ^ 13);
  assign w563[44] = |(datain[135:132] ^ 5);
  assign w563[45] = |(datain[131:128] ^ 12);
  assign w563[46] = |(datain[127:124] ^ 2);
  assign w563[47] = |(datain[123:120] ^ 14);
  assign w563[48] = |(datain[119:116] ^ 9);
  assign w563[49] = |(datain[115:112] ^ 0);
  assign w563[50] = |(datain[111:108] ^ 11);
  assign w563[51] = |(datain[107:104] ^ 4);
  assign w563[52] = |(datain[103:100] ^ 0);
  assign w563[53] = |(datain[99:96] ^ 0);
  assign w563[54] = |(datain[95:92] ^ 2);
  assign w563[55] = |(datain[91:88] ^ 14);
  assign w563[56] = |(datain[87:84] ^ 8);
  assign w563[57] = |(datain[83:80] ^ 10);
  assign w563[58] = |(datain[79:76] ^ 0);
  assign w563[59] = |(datain[75:72] ^ 7);
  assign w563[60] = |(datain[71:68] ^ 3);
  assign w563[61] = |(datain[67:64] ^ 2);
  assign w563[62] = |(datain[63:60] ^ 12);
  assign w563[63] = |(datain[59:56] ^ 4);
  assign w563[64] = |(datain[55:52] ^ 2);
  assign w563[65] = |(datain[51:48] ^ 14);
  assign w563[66] = |(datain[47:44] ^ 8);
  assign w563[67] = |(datain[43:40] ^ 8);
  assign w563[68] = |(datain[39:36] ^ 0);
  assign w563[69] = |(datain[35:32] ^ 7);
  assign w563[70] = |(datain[31:28] ^ 14);
  assign w563[71] = |(datain[27:24] ^ 8);
  assign w563[72] = |(datain[23:20] ^ 0);
  assign w563[73] = |(datain[19:16] ^ 14);
  assign w563[74] = |(datain[15:12] ^ 0);
  assign w563[75] = |(datain[11:8] ^ 0);
  assign comp[563] = ~(|w563);
  wire [32-1:0] w564;
  assign w564[0] = |(datain[311:308] ^ 0);
  assign w564[1] = |(datain[307:304] ^ 1);
  assign w564[2] = |(datain[303:300] ^ 8);
  assign w564[3] = |(datain[299:296] ^ 12);
  assign w564[4] = |(datain[295:292] ^ 12);
  assign w564[5] = |(datain[291:288] ^ 11);
  assign w564[6] = |(datain[287:284] ^ 14);
  assign w564[7] = |(datain[283:280] ^ 10);
  assign w564[8] = |(datain[279:276] ^ 0);
  assign w564[9] = |(datain[275:272] ^ 0);
  assign w564[10] = |(datain[271:268] ^ 0);
  assign w564[11] = |(datain[267:264] ^ 0);
  assign w564[12] = |(datain[263:260] ^ 0);
  assign w564[13] = |(datain[259:256] ^ 0);
  assign w564[14] = |(datain[255:252] ^ 0);
  assign w564[15] = |(datain[251:248] ^ 0);
  assign w564[16] = |(datain[247:244] ^ 8);
  assign w564[17] = |(datain[243:240] ^ 11);
  assign w564[18] = |(datain[239:236] ^ 12);
  assign w564[19] = |(datain[235:232] ^ 8);
  assign w564[20] = |(datain[231:228] ^ 8);
  assign w564[21] = |(datain[227:224] ^ 14);
  assign w564[22] = |(datain[223:220] ^ 13);
  assign w564[23] = |(datain[219:216] ^ 11);
  assign w564[24] = |(datain[215:212] ^ 11);
  assign w564[25] = |(datain[211:208] ^ 14);
  assign w564[26] = |(datain[207:204] ^ 0);
  assign w564[27] = |(datain[203:200] ^ 0);
  assign w564[28] = |(datain[199:196] ^ 0);
  assign w564[29] = |(datain[195:192] ^ 1);
  assign w564[30] = |(datain[191:188] ^ 11);
  assign w564[31] = |(datain[187:184] ^ 15);
  assign comp[564] = ~(|w564);
  wire [74-1:0] w565;
  assign w565[0] = |(datain[311:308] ^ 9);
  assign w565[1] = |(datain[307:304] ^ 14);
  assign w565[2] = |(datain[303:300] ^ 0);
  assign w565[3] = |(datain[299:296] ^ 1);
  assign w565[4] = |(datain[295:292] ^ 3);
  assign w565[5] = |(datain[291:288] ^ 9);
  assign w565[6] = |(datain[287:284] ^ 0);
  assign w565[7] = |(datain[283:280] ^ 6);
  assign w565[8] = |(datain[279:276] ^ 9);
  assign w565[9] = |(datain[275:272] ^ 12);
  assign w565[10] = |(datain[271:268] ^ 0);
  assign w565[11] = |(datain[267:264] ^ 1);
  assign w565[12] = |(datain[263:260] ^ 7);
  assign w565[13] = |(datain[259:256] ^ 4);
  assign w565[14] = |(datain[255:252] ^ 3);
  assign w565[15] = |(datain[251:248] ^ 1);
  assign w565[16] = |(datain[247:244] ^ 0);
  assign w565[17] = |(datain[243:240] ^ 5);
  assign w565[18] = |(datain[239:236] ^ 9);
  assign w565[19] = |(datain[235:232] ^ 11);
  assign w565[20] = |(datain[231:228] ^ 0);
  assign w565[21] = |(datain[227:224] ^ 1);
  assign w565[22] = |(datain[223:220] ^ 10);
  assign w565[23] = |(datain[219:216] ^ 3);
  assign w565[24] = |(datain[215:212] ^ 9);
  assign w565[25] = |(datain[211:208] ^ 9);
  assign w565[26] = |(datain[207:204] ^ 0);
  assign w565[27] = |(datain[203:200] ^ 1);
  assign w565[28] = |(datain[199:196] ^ 11);
  assign w565[29] = |(datain[195:192] ^ 8);
  assign w565[30] = |(datain[191:188] ^ 0);
  assign w565[31] = |(datain[187:184] ^ 0);
  assign w565[32] = |(datain[183:180] ^ 4);
  assign w565[33] = |(datain[179:176] ^ 2);
  assign w565[34] = |(datain[175:172] ^ 14);
  assign w565[35] = |(datain[171:168] ^ 8);
  assign w565[36] = |(datain[167:164] ^ 3);
  assign w565[37] = |(datain[163:160] ^ 10);
  assign w565[38] = |(datain[159:156] ^ 0);
  assign w565[39] = |(datain[155:152] ^ 0);
  assign w565[40] = |(datain[151:148] ^ 11);
  assign w565[41] = |(datain[147:144] ^ 8);
  assign w565[42] = |(datain[143:140] ^ 0);
  assign w565[43] = |(datain[139:136] ^ 0);
  assign w565[44] = |(datain[135:132] ^ 5);
  assign w565[45] = |(datain[131:128] ^ 7);
  assign w565[46] = |(datain[127:124] ^ 12);
  assign w565[47] = |(datain[123:120] ^ 13);
  assign w565[48] = |(datain[119:116] ^ 2);
  assign w565[49] = |(datain[115:112] ^ 1);
  assign w565[50] = |(datain[111:108] ^ 5);
  assign w565[51] = |(datain[107:104] ^ 2);
  assign w565[52] = |(datain[103:100] ^ 5);
  assign w565[53] = |(datain[99:96] ^ 1);
  assign w565[54] = |(datain[95:92] ^ 11);
  assign w565[55] = |(datain[91:88] ^ 9);
  assign w565[56] = |(datain[87:84] ^ 0);
  assign w565[57] = |(datain[83:80] ^ 3);
  assign w565[58] = |(datain[79:76] ^ 0);
  assign w565[59] = |(datain[75:72] ^ 0);
  assign w565[60] = |(datain[71:68] ^ 11);
  assign w565[61] = |(datain[67:64] ^ 4);
  assign w565[62] = |(datain[63:60] ^ 4);
  assign w565[63] = |(datain[59:56] ^ 0);
  assign w565[64] = |(datain[55:52] ^ 11);
  assign w565[65] = |(datain[51:48] ^ 10);
  assign w565[66] = |(datain[47:44] ^ 9);
  assign w565[67] = |(datain[43:40] ^ 8);
  assign w565[68] = |(datain[39:36] ^ 0);
  assign w565[69] = |(datain[35:32] ^ 1);
  assign w565[70] = |(datain[31:28] ^ 12);
  assign w565[71] = |(datain[27:24] ^ 13);
  assign w565[72] = |(datain[23:20] ^ 2);
  assign w565[73] = |(datain[19:16] ^ 1);
  assign comp[565] = ~(|w565);
  wire [74-1:0] w566;
  assign w566[0] = |(datain[311:308] ^ 8);
  assign w566[1] = |(datain[307:304] ^ 11);
  assign w566[2] = |(datain[303:300] ^ 14);
  assign w566[3] = |(datain[299:296] ^ 6);
  assign w566[4] = |(datain[295:292] ^ 8);
  assign w566[5] = |(datain[291:288] ^ 11);
  assign w566[6] = |(datain[287:284] ^ 1);
  assign w566[7] = |(datain[283:280] ^ 14);
  assign w566[8] = |(datain[279:276] ^ 1);
  assign w566[9] = |(datain[275:272] ^ 3);
  assign w566[10] = |(datain[271:268] ^ 0);
  assign w566[11] = |(datain[267:264] ^ 4);
  assign w566[12] = |(datain[263:260] ^ 8);
  assign w566[13] = |(datain[259:256] ^ 3);
  assign w566[14] = |(datain[255:252] ^ 14);
  assign w566[15] = |(datain[251:248] ^ 11);
  assign w566[16] = |(datain[247:244] ^ 0);
  assign w566[17] = |(datain[243:240] ^ 3);
  assign w566[18] = |(datain[239:236] ^ 11);
  assign w566[19] = |(datain[235:232] ^ 1);
  assign w566[20] = |(datain[231:228] ^ 0);
  assign w566[21] = |(datain[227:224] ^ 6);
  assign w566[22] = |(datain[223:220] ^ 8);
  assign w566[23] = |(datain[219:216] ^ 9);
  assign w566[24] = |(datain[215:212] ^ 1);
  assign w566[25] = |(datain[211:208] ^ 14);
  assign w566[26] = |(datain[207:204] ^ 1);
  assign w566[27] = |(datain[203:200] ^ 3);
  assign w566[28] = |(datain[199:196] ^ 0);
  assign w566[29] = |(datain[195:192] ^ 4);
  assign w566[30] = |(datain[191:188] ^ 13);
  assign w566[31] = |(datain[187:184] ^ 3);
  assign w566[32] = |(datain[183:180] ^ 14);
  assign w566[33] = |(datain[179:176] ^ 3);
  assign w566[34] = |(datain[175:172] ^ 8);
  assign w566[35] = |(datain[171:168] ^ 3);
  assign w566[36] = |(datain[167:164] ^ 14);
  assign w566[37] = |(datain[163:160] ^ 11);
  assign w566[38] = |(datain[159:156] ^ 1);
  assign w566[39] = |(datain[155:152] ^ 0);
  assign w566[40] = |(datain[151:148] ^ 8);
  assign w566[41] = |(datain[147:144] ^ 14);
  assign w566[42] = |(datain[143:140] ^ 12);
  assign w566[43] = |(datain[139:136] ^ 3);
  assign w566[44] = |(datain[135:132] ^ 11);
  assign w566[45] = |(datain[131:128] ^ 9);
  assign w566[46] = |(datain[127:124] ^ 0);
  assign w566[47] = |(datain[123:120] ^ 0);
  assign w566[48] = |(datain[119:116] ^ 0);
  assign w566[49] = |(datain[115:112] ^ 1);
  assign w566[50] = |(datain[111:108] ^ 8);
  assign w566[51] = |(datain[107:104] ^ 11);
  assign w566[52] = |(datain[103:100] ^ 15);
  assign w566[53] = |(datain[99:96] ^ 9);
  assign w566[54] = |(datain[95:92] ^ 15);
  assign w566[55] = |(datain[91:88] ^ 3);
  assign w566[56] = |(datain[87:84] ^ 10);
  assign w566[57] = |(datain[83:80] ^ 5);
  assign w566[58] = |(datain[79:76] ^ 0);
  assign w566[59] = |(datain[75:72] ^ 6);
  assign w566[60] = |(datain[71:68] ^ 14);
  assign w566[61] = |(datain[67:64] ^ 8);
  assign w566[62] = |(datain[63:60] ^ 0);
  assign w566[63] = |(datain[59:56] ^ 0);
  assign w566[64] = |(datain[55:52] ^ 0);
  assign w566[65] = |(datain[51:48] ^ 0);
  assign w566[66] = |(datain[47:44] ^ 5);
  assign w566[67] = |(datain[43:40] ^ 9);
  assign w566[68] = |(datain[39:36] ^ 8);
  assign w566[69] = |(datain[35:32] ^ 1);
  assign w566[70] = |(datain[31:28] ^ 14);
  assign w566[71] = |(datain[27:24] ^ 9);
  assign w566[72] = |(datain[23:20] ^ 15);
  assign w566[73] = |(datain[19:16] ^ 9);
  assign comp[566] = ~(|w566);
  wire [40-1:0] w567;
  assign w567[0] = |(datain[311:308] ^ 0);
  assign w567[1] = |(datain[307:304] ^ 3);
  assign w567[2] = |(datain[303:300] ^ 1);
  assign w567[3] = |(datain[299:296] ^ 14);
  assign w567[4] = |(datain[295:292] ^ 0);
  assign w567[5] = |(datain[291:288] ^ 6);
  assign w567[6] = |(datain[287:284] ^ 3);
  assign w567[7] = |(datain[283:280] ^ 3);
  assign w567[8] = |(datain[279:276] ^ 12);
  assign w567[9] = |(datain[275:272] ^ 0);
  assign w567[10] = |(datain[271:268] ^ 5);
  assign w567[11] = |(datain[267:264] ^ 0);
  assign w567[12] = |(datain[263:260] ^ 1);
  assign w567[13] = |(datain[259:256] ^ 15);
  assign w567[14] = |(datain[255:252] ^ 11);
  assign w567[15] = |(datain[251:248] ^ 14);
  assign w567[16] = |(datain[247:244] ^ 8);
  assign w567[17] = |(datain[243:240] ^ 4);
  assign w567[18] = |(datain[239:236] ^ 0);
  assign w567[19] = |(datain[235:232] ^ 0);
  assign w567[20] = |(datain[231:228] ^ 8);
  assign w567[21] = |(datain[227:224] ^ 11);
  assign w567[22] = |(datain[223:220] ^ 4);
  assign w567[23] = |(datain[219:216] ^ 4);
  assign w567[24] = |(datain[215:212] ^ 0);
  assign w567[25] = |(datain[211:208] ^ 2);
  assign w567[26] = |(datain[207:204] ^ 8);
  assign w567[27] = |(datain[203:200] ^ 14);
  assign w567[28] = |(datain[199:196] ^ 12);
  assign w567[29] = |(datain[195:192] ^ 0);
  assign w567[30] = |(datain[191:188] ^ 8);
  assign w567[31] = |(datain[187:184] ^ 11);
  assign w567[32] = |(datain[183:180] ^ 3);
  assign w567[33] = |(datain[179:176] ^ 12);
  assign w567[34] = |(datain[175:172] ^ 2);
  assign w567[35] = |(datain[171:168] ^ 6);
  assign w567[36] = |(datain[167:164] ^ 8);
  assign w567[37] = |(datain[163:160] ^ 1);
  assign w567[38] = |(datain[159:156] ^ 7);
  assign w567[39] = |(datain[155:152] ^ 13);
  assign comp[567] = ~(|w567);
  wire [74-1:0] w568;
  assign w568[0] = |(datain[311:308] ^ 8);
  assign w568[1] = |(datain[307:304] ^ 12);
  assign w568[2] = |(datain[303:300] ^ 12);
  assign w568[3] = |(datain[299:296] ^ 8);
  assign w568[4] = |(datain[295:292] ^ 8);
  assign w568[5] = |(datain[291:288] ^ 14);
  assign w568[6] = |(datain[287:284] ^ 13);
  assign w568[7] = |(datain[283:280] ^ 8);
  assign w568[8] = |(datain[279:276] ^ 8);
  assign w568[9] = |(datain[275:272] ^ 12);
  assign w568[10] = |(datain[271:268] ^ 0);
  assign w568[11] = |(datain[267:264] ^ 6);
  assign w568[12] = |(datain[263:260] ^ 7);
  assign w568[13] = |(datain[259:256] ^ 3);
  assign w568[14] = |(datain[255:252] ^ 0);
  assign w568[15] = |(datain[251:248] ^ 9);
  assign w568[16] = |(datain[247:244] ^ 8);
  assign w568[17] = |(datain[243:240] ^ 12);
  assign w568[18] = |(datain[239:236] ^ 1);
  assign w568[19] = |(datain[235:232] ^ 6);
  assign w568[20] = |(datain[231:228] ^ 7);
  assign w568[21] = |(datain[227:224] ^ 1);
  assign w568[22] = |(datain[223:220] ^ 0);
  assign w568[23] = |(datain[219:216] ^ 9);
  assign w568[24] = |(datain[215:212] ^ 8);
  assign w568[25] = |(datain[211:208] ^ 9);
  assign w568[26] = |(datain[207:204] ^ 2);
  assign w568[27] = |(datain[203:200] ^ 6);
  assign w568[28] = |(datain[199:196] ^ 6);
  assign w568[29] = |(datain[195:192] ^ 15);
  assign w568[30] = |(datain[191:188] ^ 0);
  assign w568[31] = |(datain[187:184] ^ 9);
  assign w568[32] = |(datain[183:180] ^ 8);
  assign w568[33] = |(datain[179:176] ^ 14);
  assign w568[34] = |(datain[175:172] ^ 13);
  assign w568[35] = |(datain[171:168] ^ 0);
  assign w568[36] = |(datain[167:164] ^ 11);
  assign w568[37] = |(datain[163:160] ^ 12);
  assign w568[38] = |(datain[159:156] ^ 5);
  assign w568[39] = |(datain[155:152] ^ 6);
  assign w568[40] = |(datain[151:148] ^ 0);
  assign w568[41] = |(datain[147:144] ^ 10);
  assign w568[42] = |(datain[143:140] ^ 15);
  assign w568[43] = |(datain[139:136] ^ 11);
  assign w568[44] = |(datain[135:132] ^ 10);
  assign w568[45] = |(datain[131:128] ^ 1);
  assign w568[46] = |(datain[127:124] ^ 6);
  assign w568[47] = |(datain[123:120] ^ 1);
  assign w568[48] = |(datain[119:116] ^ 0);
  assign w568[49] = |(datain[115:112] ^ 9);
  assign w568[50] = |(datain[111:108] ^ 11);
  assign w568[51] = |(datain[107:104] ^ 14);
  assign w568[52] = |(datain[103:100] ^ 4);
  assign w568[53] = |(datain[99:96] ^ 6);
  assign w568[54] = |(datain[95:92] ^ 0);
  assign w568[55] = |(datain[91:88] ^ 1);
  assign w568[56] = |(datain[87:84] ^ 11);
  assign w568[57] = |(datain[83:80] ^ 9);
  assign w568[58] = |(datain[79:76] ^ 3);
  assign w568[59] = |(datain[75:72] ^ 15);
  assign w568[60] = |(datain[71:68] ^ 0);
  assign w568[61] = |(datain[67:64] ^ 9);
  assign w568[62] = |(datain[63:60] ^ 12);
  assign w568[63] = |(datain[59:56] ^ 6);
  assign w568[64] = |(datain[55:52] ^ 0);
  assign w568[65] = |(datain[51:48] ^ 6);
  assign w568[66] = |(datain[47:44] ^ 0);
  assign w568[67] = |(datain[43:40] ^ 15);
  assign w568[68] = |(datain[39:36] ^ 0);
  assign w568[69] = |(datain[35:32] ^ 1);
  assign w568[70] = |(datain[31:28] ^ 3);
  assign w568[71] = |(datain[27:24] ^ 0);
  assign w568[72] = |(datain[23:20] ^ 14);
  assign w568[73] = |(datain[19:16] ^ 8);
  assign comp[568] = ~(|w568);
  wire [44-1:0] w569;
  assign w569[0] = |(datain[311:308] ^ 4);
  assign w569[1] = |(datain[307:304] ^ 4);
  assign w569[2] = |(datain[303:300] ^ 7);
  assign w569[3] = |(datain[299:296] ^ 4);
  assign w569[4] = |(datain[295:292] ^ 14);
  assign w569[5] = |(datain[291:288] ^ 4);
  assign w569[6] = |(datain[287:284] ^ 5);
  assign w569[7] = |(datain[283:280] ^ 0);
  assign w569[8] = |(datain[279:276] ^ 5);
  assign w569[9] = |(datain[275:272] ^ 3);
  assign w569[10] = |(datain[271:268] ^ 5);
  assign w569[11] = |(datain[267:264] ^ 1);
  assign w569[12] = |(datain[263:260] ^ 0);
  assign w569[13] = |(datain[259:256] ^ 6);
  assign w569[14] = |(datain[255:252] ^ 5);
  assign w569[15] = |(datain[251:248] ^ 6);
  assign w569[16] = |(datain[247:244] ^ 5);
  assign w569[17] = |(datain[243:240] ^ 7);
  assign w569[18] = |(datain[239:236] ^ 5);
  assign w569[19] = |(datain[235:232] ^ 2);
  assign w569[20] = |(datain[231:228] ^ 1);
  assign w569[21] = |(datain[227:224] ^ 14);
  assign w569[22] = |(datain[223:220] ^ 5);
  assign w569[23] = |(datain[219:216] ^ 5);
  assign w569[24] = |(datain[215:212] ^ 8);
  assign w569[25] = |(datain[211:208] ^ 0);
  assign w569[26] = |(datain[207:204] ^ 15);
  assign w569[27] = |(datain[203:200] ^ 12);
  assign w569[28] = |(datain[199:196] ^ 6);
  assign w569[29] = |(datain[195:192] ^ 12);
  assign w569[30] = |(datain[191:188] ^ 7);
  assign w569[31] = |(datain[187:184] ^ 4);
  assign w569[32] = |(datain[183:180] ^ 1);
  assign w569[33] = |(datain[179:176] ^ 6);
  assign w569[34] = |(datain[175:172] ^ 3);
  assign w569[35] = |(datain[171:168] ^ 13);
  assign w569[36] = |(datain[167:164] ^ 0);
  assign w569[37] = |(datain[163:160] ^ 0);
  assign w569[38] = |(datain[159:156] ^ 4);
  assign w569[39] = |(datain[155:152] ^ 11);
  assign w569[40] = |(datain[151:148] ^ 7);
  assign w569[41] = |(datain[147:144] ^ 4);
  assign w569[42] = |(datain[143:140] ^ 0);
  assign w569[43] = |(datain[139:136] ^ 15);
  assign comp[569] = ~(|w569);
  wire [46-1:0] w570;
  assign w570[0] = |(datain[311:308] ^ 8);
  assign w570[1] = |(datain[307:304] ^ 14);
  assign w570[2] = |(datain[303:300] ^ 13);
  assign w570[3] = |(datain[299:296] ^ 8);
  assign w570[4] = |(datain[295:292] ^ 8);
  assign w570[5] = |(datain[291:288] ^ 11);
  assign w570[6] = |(datain[287:284] ^ 1);
  assign w570[7] = |(datain[283:280] ^ 14);
  assign w570[8] = |(datain[279:276] ^ 0);
  assign w570[9] = |(datain[275:272] ^ 3);
  assign w570[10] = |(datain[271:268] ^ 0);
  assign w570[11] = |(datain[267:264] ^ 0);
  assign w570[12] = |(datain[263:260] ^ 3);
  assign w570[13] = |(datain[259:256] ^ 3);
  assign w570[14] = |(datain[255:252] ^ 15);
  assign w570[15] = |(datain[251:248] ^ 15);
  assign w570[16] = |(datain[247:244] ^ 11);
  assign w570[17] = |(datain[243:240] ^ 9);
  assign w570[18] = |(datain[239:236] ^ 3);
  assign w570[19] = |(datain[235:232] ^ 1);
  assign w570[20] = |(datain[231:228] ^ 0);
  assign w570[21] = |(datain[227:224] ^ 3);
  assign w570[22] = |(datain[223:220] ^ 11);
  assign w570[23] = |(datain[219:216] ^ 8);
  assign w570[24] = |(datain[215:212] ^ 10);
  assign w570[25] = |(datain[211:208] ^ 9);
  assign w570[26] = |(datain[207:204] ^ 4);
  assign w570[27] = |(datain[203:200] ^ 4);
  assign w570[28] = |(datain[199:196] ^ 12);
  assign w570[29] = |(datain[195:192] ^ 13);
  assign w570[30] = |(datain[191:188] ^ 2);
  assign w570[31] = |(datain[187:184] ^ 1);
  assign w570[32] = |(datain[183:180] ^ 7);
  assign w570[33] = |(datain[179:176] ^ 3);
  assign w570[34] = |(datain[175:172] ^ 7);
  assign w570[35] = |(datain[171:168] ^ 12);
  assign w570[36] = |(datain[167:164] ^ 11);
  assign w570[37] = |(datain[163:160] ^ 8);
  assign w570[38] = |(datain[159:156] ^ 4);
  assign w570[39] = |(datain[155:152] ^ 4);
  assign w570[40] = |(datain[151:148] ^ 0);
  assign w570[41] = |(datain[147:144] ^ 0);
  assign w570[42] = |(datain[143:140] ^ 8);
  assign w570[43] = |(datain[139:136] ^ 5);
  assign w570[44] = |(datain[135:132] ^ 14);
  assign w570[45] = |(datain[131:128] ^ 13);
  assign comp[570] = ~(|w570);
  wire [74-1:0] w571;
  assign w571[0] = |(datain[311:308] ^ 10);
  assign w571[1] = |(datain[307:304] ^ 3);
  assign w571[2] = |(datain[303:300] ^ 0);
  assign w571[3] = |(datain[299:296] ^ 12);
  assign w571[4] = |(datain[295:292] ^ 7);
  assign w571[5] = |(datain[291:288] ^ 13);
  assign w571[6] = |(datain[287:284] ^ 10);
  assign w571[7] = |(datain[283:280] ^ 1);
  assign w571[8] = |(datain[279:276] ^ 4);
  assign w571[9] = |(datain[275:272] ^ 14);
  assign w571[10] = |(datain[271:268] ^ 0);
  assign w571[11] = |(datain[267:264] ^ 0);
  assign w571[12] = |(datain[263:260] ^ 10);
  assign w571[13] = |(datain[259:256] ^ 3);
  assign w571[14] = |(datain[255:252] ^ 0);
  assign w571[15] = |(datain[251:248] ^ 14);
  assign w571[16] = |(datain[247:244] ^ 7);
  assign w571[17] = |(datain[243:240] ^ 13);
  assign w571[18] = |(datain[239:236] ^ 11);
  assign w571[19] = |(datain[235:232] ^ 11);
  assign w571[20] = |(datain[231:228] ^ 4);
  assign w571[21] = |(datain[227:224] ^ 12);
  assign w571[22] = |(datain[223:220] ^ 0);
  assign w571[23] = |(datain[219:216] ^ 0);
  assign w571[24] = |(datain[215:212] ^ 8);
  assign w571[25] = |(datain[211:208] ^ 11);
  assign w571[26] = |(datain[207:204] ^ 8);
  assign w571[27] = |(datain[203:200] ^ 7);
  assign w571[28] = |(datain[199:196] ^ 12);
  assign w571[29] = |(datain[195:192] ^ 7);
  assign w571[30] = |(datain[191:188] ^ 0);
  assign w571[31] = |(datain[187:184] ^ 3);
  assign w571[32] = |(datain[183:180] ^ 4);
  assign w571[33] = |(datain[179:176] ^ 8);
  assign w571[34] = |(datain[175:172] ^ 8);
  assign w571[35] = |(datain[171:168] ^ 9);
  assign w571[36] = |(datain[167:164] ^ 8);
  assign w571[37] = |(datain[163:160] ^ 7);
  assign w571[38] = |(datain[159:156] ^ 12);
  assign w571[39] = |(datain[155:152] ^ 7);
  assign w571[40] = |(datain[151:148] ^ 0);
  assign w571[41] = |(datain[147:144] ^ 3);
  assign w571[42] = |(datain[143:140] ^ 12);
  assign w571[43] = |(datain[139:136] ^ 1);
  assign w571[44] = |(datain[135:132] ^ 14);
  assign w571[45] = |(datain[131:128] ^ 0);
  assign w571[46] = |(datain[127:124] ^ 0);
  assign w571[47] = |(datain[123:120] ^ 6);
  assign w571[48] = |(datain[119:116] ^ 8);
  assign w571[49] = |(datain[115:112] ^ 9);
  assign w571[50] = |(datain[111:108] ^ 4);
  assign w571[51] = |(datain[107:104] ^ 7);
  assign w571[52] = |(datain[103:100] ^ 0);
  assign w571[53] = |(datain[99:96] ^ 2);
  assign w571[54] = |(datain[95:92] ^ 12);
  assign w571[55] = |(datain[91:88] ^ 7);
  assign w571[56] = |(datain[87:84] ^ 0);
  assign w571[57] = |(datain[83:80] ^ 7);
  assign w571[58] = |(datain[79:76] ^ 7);
  assign w571[59] = |(datain[75:72] ^ 3);
  assign w571[60] = |(datain[71:68] ^ 0);
  assign w571[61] = |(datain[67:64] ^ 1);
  assign w571[62] = |(datain[63:60] ^ 10);
  assign w571[63] = |(datain[59:56] ^ 3);
  assign w571[64] = |(datain[55:52] ^ 2);
  assign w571[65] = |(datain[51:48] ^ 6);
  assign w571[66] = |(datain[47:44] ^ 0);
  assign w571[67] = |(datain[43:40] ^ 0);
  assign w571[68] = |(datain[39:36] ^ 12);
  assign w571[69] = |(datain[35:32] ^ 7);
  assign w571[70] = |(datain[31:28] ^ 0);
  assign w571[71] = |(datain[27:24] ^ 6);
  assign w571[72] = |(datain[23:20] ^ 2);
  assign w571[73] = |(datain[19:16] ^ 4);
  assign comp[571] = ~(|w571);
  wire [46-1:0] w572;
  assign w572[0] = |(datain[311:308] ^ 0);
  assign w572[1] = |(datain[307:304] ^ 2);
  assign w572[2] = |(datain[303:300] ^ 0);
  assign w572[3] = |(datain[299:296] ^ 0);
  assign w572[4] = |(datain[295:292] ^ 14);
  assign w572[5] = |(datain[291:288] ^ 11);
  assign w572[6] = |(datain[287:284] ^ 2);
  assign w572[7] = |(datain[283:280] ^ 1);
  assign w572[8] = |(datain[279:276] ^ 3);
  assign w572[9] = |(datain[275:272] ^ 14);
  assign w572[10] = |(datain[271:268] ^ 8);
  assign w572[11] = |(datain[267:264] ^ 10);
  assign w572[12] = |(datain[263:260] ^ 8);
  assign w572[13] = |(datain[259:256] ^ 6);
  assign w572[14] = |(datain[255:252] ^ 4);
  assign w572[15] = |(datain[251:248] ^ 6);
  assign w572[16] = |(datain[247:244] ^ 0);
  assign w572[17] = |(datain[243:240] ^ 7);
  assign w572[18] = |(datain[239:236] ^ 8);
  assign w572[19] = |(datain[235:232] ^ 13);
  assign w572[20] = |(datain[231:228] ^ 11);
  assign w572[21] = |(datain[227:224] ^ 6);
  assign w572[22] = |(datain[223:220] ^ 3);
  assign w572[23] = |(datain[219:216] ^ 5);
  assign w572[24] = |(datain[215:212] ^ 0);
  assign w572[25] = |(datain[211:208] ^ 1);
  assign w572[26] = |(datain[207:204] ^ 11);
  assign w572[27] = |(datain[203:200] ^ 9);
  assign w572[28] = |(datain[199:196] ^ 0);
  assign w572[29] = |(datain[195:192] ^ 15);
  assign w572[30] = |(datain[191:188] ^ 0);
  assign w572[31] = |(datain[187:184] ^ 6);
  assign w572[32] = |(datain[183:180] ^ 3);
  assign w572[33] = |(datain[179:176] ^ 0);
  assign w572[34] = |(datain[175:172] ^ 0);
  assign w572[35] = |(datain[171:168] ^ 4);
  assign w572[36] = |(datain[167:164] ^ 13);
  assign w572[37] = |(datain[163:160] ^ 2);
  assign w572[38] = |(datain[159:156] ^ 12);
  assign w572[39] = |(datain[155:152] ^ 0);
  assign w572[40] = |(datain[151:148] ^ 4);
  assign w572[41] = |(datain[147:144] ^ 6);
  assign w572[42] = |(datain[143:140] ^ 14);
  assign w572[43] = |(datain[139:136] ^ 2);
  assign w572[44] = |(datain[135:132] ^ 15);
  assign w572[45] = |(datain[131:128] ^ 9);
  assign comp[572] = ~(|w572);
  wire [46-1:0] w573;
  assign w573[0] = |(datain[311:308] ^ 0);
  assign w573[1] = |(datain[307:304] ^ 2);
  assign w573[2] = |(datain[303:300] ^ 0);
  assign w573[3] = |(datain[299:296] ^ 0);
  assign w573[4] = |(datain[295:292] ^ 14);
  assign w573[5] = |(datain[291:288] ^ 11);
  assign w573[6] = |(datain[287:284] ^ 2);
  assign w573[7] = |(datain[283:280] ^ 1);
  assign w573[8] = |(datain[279:276] ^ 3);
  assign w573[9] = |(datain[275:272] ^ 14);
  assign w573[10] = |(datain[271:268] ^ 8);
  assign w573[11] = |(datain[267:264] ^ 10);
  assign w573[12] = |(datain[263:260] ^ 8);
  assign w573[13] = |(datain[259:256] ^ 6);
  assign w573[14] = |(datain[255:252] ^ 4);
  assign w573[15] = |(datain[251:248] ^ 9);
  assign w573[16] = |(datain[247:244] ^ 0);
  assign w573[17] = |(datain[243:240] ^ 7);
  assign w573[18] = |(datain[239:236] ^ 8);
  assign w573[19] = |(datain[235:232] ^ 13);
  assign w573[20] = |(datain[231:228] ^ 11);
  assign w573[21] = |(datain[227:224] ^ 6);
  assign w573[22] = |(datain[223:220] ^ 3);
  assign w573[23] = |(datain[219:216] ^ 6);
  assign w573[24] = |(datain[215:212] ^ 0);
  assign w573[25] = |(datain[211:208] ^ 1);
  assign w573[26] = |(datain[207:204] ^ 11);
  assign w573[27] = |(datain[203:200] ^ 9);
  assign w573[28] = |(datain[199:196] ^ 1);
  assign w573[29] = |(datain[195:192] ^ 1);
  assign w573[30] = |(datain[191:188] ^ 0);
  assign w573[31] = |(datain[187:184] ^ 6);
  assign w573[32] = |(datain[183:180] ^ 3);
  assign w573[33] = |(datain[179:176] ^ 0);
  assign w573[34] = |(datain[175:172] ^ 0);
  assign w573[35] = |(datain[171:168] ^ 4);
  assign w573[36] = |(datain[167:164] ^ 13);
  assign w573[37] = |(datain[163:160] ^ 2);
  assign w573[38] = |(datain[159:156] ^ 12);
  assign w573[39] = |(datain[155:152] ^ 0);
  assign w573[40] = |(datain[151:148] ^ 4);
  assign w573[41] = |(datain[147:144] ^ 6);
  assign w573[42] = |(datain[143:140] ^ 14);
  assign w573[43] = |(datain[139:136] ^ 2);
  assign w573[44] = |(datain[135:132] ^ 15);
  assign w573[45] = |(datain[131:128] ^ 9);
  assign comp[573] = ~(|w573);
  wire [34-1:0] w574;
  assign w574[0] = |(datain[311:308] ^ 0);
  assign w574[1] = |(datain[307:304] ^ 2);
  assign w574[2] = |(datain[303:300] ^ 8);
  assign w574[3] = |(datain[299:296] ^ 13);
  assign w574[4] = |(datain[295:292] ^ 11);
  assign w574[5] = |(datain[291:288] ^ 6);
  assign w574[6] = |(datain[287:284] ^ 3);
  assign w574[7] = |(datain[283:280] ^ 10);
  assign w574[8] = |(datain[279:276] ^ 0);
  assign w574[9] = |(datain[275:272] ^ 2);
  assign w574[10] = |(datain[271:268] ^ 5);
  assign w574[11] = |(datain[267:264] ^ 2);
  assign w574[12] = |(datain[263:260] ^ 14);
  assign w574[13] = |(datain[259:256] ^ 11);
  assign w574[14] = |(datain[255:252] ^ 2);
  assign w574[15] = |(datain[251:248] ^ 9);
  assign w574[16] = |(datain[247:244] ^ 11);
  assign w574[17] = |(datain[243:240] ^ 4);
  assign w574[18] = |(datain[239:236] ^ 1);
  assign w574[19] = |(datain[235:232] ^ 10);
  assign w574[20] = |(datain[231:228] ^ 11);
  assign w574[21] = |(datain[227:224] ^ 10);
  assign w574[22] = |(datain[223:220] ^ 8);
  assign w574[23] = |(datain[219:216] ^ 0);
  assign w574[24] = |(datain[215:212] ^ 0);
  assign w574[25] = |(datain[211:208] ^ 0);
  assign w574[26] = |(datain[207:204] ^ 12);
  assign w574[27] = |(datain[203:200] ^ 13);
  assign w574[28] = |(datain[199:196] ^ 2);
  assign w574[29] = |(datain[195:192] ^ 1);
  assign w574[30] = |(datain[191:188] ^ 3);
  assign w574[31] = |(datain[187:184] ^ 3);
  assign w574[32] = |(datain[183:180] ^ 12);
  assign w574[33] = |(datain[179:176] ^ 0);
  assign comp[574] = ~(|w574);
  wire [42-1:0] w575;
  assign w575[0] = |(datain[311:308] ^ 5);
  assign w575[1] = |(datain[307:304] ^ 13);
  assign w575[2] = |(datain[303:300] ^ 8);
  assign w575[3] = |(datain[299:296] ^ 1);
  assign w575[4] = |(datain[295:292] ^ 14);
  assign w575[5] = |(datain[291:288] ^ 13);
  assign w575[6] = |(datain[287:284] ^ 0);
  assign w575[7] = |(datain[283:280] ^ 11);
  assign w575[8] = |(datain[279:276] ^ 0);
  assign w575[9] = |(datain[275:272] ^ 1);
  assign w575[10] = |(datain[271:268] ^ 11);
  assign w575[11] = |(datain[267:264] ^ 15);
  assign w575[12] = |(datain[263:260] ^ 0);
  assign w575[13] = |(datain[259:256] ^ 0);
  assign w575[14] = |(datain[255:252] ^ 0);
  assign w575[15] = |(datain[251:248] ^ 1);
  assign w575[16] = |(datain[247:244] ^ 8);
  assign w575[17] = |(datain[243:240] ^ 13);
  assign w575[18] = |(datain[239:236] ^ 11);
  assign w575[19] = |(datain[235:232] ^ 6);
  assign w575[20] = |(datain[231:228] ^ 0);
  assign w575[21] = |(datain[227:224] ^ 4);
  assign w575[22] = |(datain[223:220] ^ 0);
  assign w575[23] = |(datain[219:216] ^ 1);
  assign w575[24] = |(datain[215:212] ^ 11);
  assign w575[25] = |(datain[211:208] ^ 9);
  assign w575[26] = |(datain[207:204] ^ 0);
  assign w575[27] = |(datain[203:200] ^ 4);
  assign w575[28] = |(datain[199:196] ^ 0);
  assign w575[29] = |(datain[195:192] ^ 0);
  assign w575[30] = |(datain[191:188] ^ 15);
  assign w575[31] = |(datain[187:184] ^ 12);
  assign w575[32] = |(datain[183:180] ^ 15);
  assign w575[33] = |(datain[179:176] ^ 3);
  assign w575[34] = |(datain[175:172] ^ 10);
  assign w575[35] = |(datain[171:168] ^ 4);
  assign w575[36] = |(datain[167:164] ^ 11);
  assign w575[37] = |(datain[163:160] ^ 4);
  assign w575[38] = |(datain[159:156] ^ 1);
  assign w575[39] = |(datain[155:152] ^ 10);
  assign w575[40] = |(datain[151:148] ^ 8);
  assign w575[41] = |(datain[147:144] ^ 13);
  assign comp[575] = ~(|w575);
  wire [32-1:0] w576;
  assign w576[0] = |(datain[311:308] ^ 8);
  assign w576[1] = |(datain[307:304] ^ 13);
  assign w576[2] = |(datain[303:300] ^ 11);
  assign w576[3] = |(datain[299:296] ^ 6);
  assign w576[4] = |(datain[295:292] ^ 3);
  assign w576[5] = |(datain[291:288] ^ 10);
  assign w576[6] = |(datain[287:284] ^ 0);
  assign w576[7] = |(datain[283:280] ^ 2);
  assign w576[8] = |(datain[279:276] ^ 5);
  assign w576[9] = |(datain[275:272] ^ 2);
  assign w576[10] = |(datain[271:268] ^ 14);
  assign w576[11] = |(datain[267:264] ^ 11);
  assign w576[12] = |(datain[263:260] ^ 2);
  assign w576[13] = |(datain[259:256] ^ 9);
  assign w576[14] = |(datain[255:252] ^ 11);
  assign w576[15] = |(datain[251:248] ^ 4);
  assign w576[16] = |(datain[247:244] ^ 1);
  assign w576[17] = |(datain[243:240] ^ 10);
  assign w576[18] = |(datain[239:236] ^ 11);
  assign w576[19] = |(datain[235:232] ^ 10);
  assign w576[20] = |(datain[231:228] ^ 8);
  assign w576[21] = |(datain[227:224] ^ 0);
  assign w576[22] = |(datain[223:220] ^ 0);
  assign w576[23] = |(datain[219:216] ^ 0);
  assign w576[24] = |(datain[215:212] ^ 12);
  assign w576[25] = |(datain[211:208] ^ 13);
  assign w576[26] = |(datain[207:204] ^ 2);
  assign w576[27] = |(datain[203:200] ^ 1);
  assign w576[28] = |(datain[199:196] ^ 3);
  assign w576[29] = |(datain[195:192] ^ 3);
  assign w576[30] = |(datain[191:188] ^ 12);
  assign w576[31] = |(datain[187:184] ^ 0);
  assign comp[576] = ~(|w576);
  wire [42-1:0] w577;
  assign w577[0] = |(datain[311:308] ^ 0);
  assign w577[1] = |(datain[307:304] ^ 1);
  assign w577[2] = |(datain[303:300] ^ 11);
  assign w577[3] = |(datain[299:296] ^ 9);
  assign w577[4] = |(datain[295:292] ^ 2);
  assign w577[5] = |(datain[291:288] ^ 10);
  assign w577[6] = |(datain[287:284] ^ 0);
  assign w577[7] = |(datain[283:280] ^ 1);
  assign w577[8] = |(datain[279:276] ^ 11);
  assign w577[9] = |(datain[275:272] ^ 4);
  assign w577[10] = |(datain[271:268] ^ 4);
  assign w577[11] = |(datain[267:264] ^ 0);
  assign w577[12] = |(datain[263:260] ^ 12);
  assign w577[13] = |(datain[259:256] ^ 13);
  assign w577[14] = |(datain[255:252] ^ 2);
  assign w577[15] = |(datain[251:248] ^ 1);
  assign w577[16] = |(datain[247:244] ^ 11);
  assign w577[17] = |(datain[243:240] ^ 8);
  assign w577[18] = |(datain[239:236] ^ 0);
  assign w577[19] = |(datain[235:232] ^ 0);
  assign w577[20] = |(datain[231:228] ^ 4);
  assign w577[21] = |(datain[227:224] ^ 2);
  assign w577[22] = |(datain[223:220] ^ 9);
  assign w577[23] = |(datain[219:216] ^ 9);
  assign w577[24] = |(datain[215:212] ^ 3);
  assign w577[25] = |(datain[211:208] ^ 3);
  assign w577[26] = |(datain[207:204] ^ 12);
  assign w577[27] = |(datain[203:200] ^ 9);
  assign w577[28] = |(datain[199:196] ^ 12);
  assign w577[29] = |(datain[195:192] ^ 13);
  assign w577[30] = |(datain[191:188] ^ 2);
  assign w577[31] = |(datain[187:184] ^ 1);
  assign w577[32] = |(datain[183:180] ^ 8);
  assign w577[33] = |(datain[179:176] ^ 11);
  assign w577[34] = |(datain[175:172] ^ 8);
  assign w577[35] = |(datain[171:168] ^ 6);
  assign w577[36] = |(datain[167:164] ^ 3);
  assign w577[37] = |(datain[163:160] ^ 13);
  assign w577[38] = |(datain[159:156] ^ 0);
  assign w577[39] = |(datain[155:152] ^ 2);
  assign w577[40] = |(datain[151:148] ^ 4);
  assign w577[41] = |(datain[147:144] ^ 0);
  assign comp[577] = ~(|w577);
  wire [60-1:0] w578;
  assign w578[0] = |(datain[311:308] ^ 9);
  assign w578[1] = |(datain[307:304] ^ 0);
  assign w578[2] = |(datain[303:300] ^ 9);
  assign w578[3] = |(datain[299:296] ^ 0);
  assign w578[4] = |(datain[295:292] ^ 12);
  assign w578[5] = |(datain[291:288] ^ 13);
  assign w578[6] = |(datain[287:284] ^ 2);
  assign w578[7] = |(datain[283:280] ^ 0);
  assign w578[8] = |(datain[279:276] ^ 9);
  assign w578[9] = |(datain[275:272] ^ 0);
  assign w578[10] = |(datain[271:268] ^ 0);
  assign w578[11] = |(datain[267:264] ^ 1);
  assign w578[12] = |(datain[263:260] ^ 14);
  assign w578[13] = |(datain[259:256] ^ 8);
  assign w578[14] = |(datain[255:252] ^ 0);
  assign w578[15] = |(datain[251:248] ^ 0);
  assign w578[16] = |(datain[247:244] ^ 0);
  assign w578[17] = |(datain[243:240] ^ 0);
  assign w578[18] = |(datain[239:236] ^ 5);
  assign w578[19] = |(datain[235:232] ^ 13);
  assign w578[20] = |(datain[231:228] ^ 8);
  assign w578[21] = |(datain[227:224] ^ 1);
  assign w578[22] = |(datain[223:220] ^ 14);
  assign w578[23] = |(datain[219:216] ^ 13);
  assign w578[24] = |(datain[215:212] ^ 0);
  assign w578[25] = |(datain[211:208] ^ 11);
  assign w578[26] = |(datain[207:204] ^ 0);
  assign w578[27] = |(datain[203:200] ^ 1);
  assign w578[28] = |(datain[199:196] ^ 11);
  assign w578[29] = |(datain[195:192] ^ 15);
  assign w578[30] = |(datain[191:188] ^ 0);
  assign w578[31] = |(datain[187:184] ^ 0);
  assign w578[32] = |(datain[183:180] ^ 0);
  assign w578[33] = |(datain[179:176] ^ 1);
  assign w578[34] = |(datain[175:172] ^ 8);
  assign w578[35] = |(datain[171:168] ^ 13);
  assign w578[36] = |(datain[167:164] ^ 11);
  assign w578[37] = |(datain[163:160] ^ 6);
  assign w578[38] = |(datain[159:156] ^ 0);
  assign w578[39] = |(datain[155:152] ^ 4);
  assign w578[40] = |(datain[151:148] ^ 0);
  assign w578[41] = |(datain[147:144] ^ 1);
  assign w578[42] = |(datain[143:140] ^ 11);
  assign w578[43] = |(datain[139:136] ^ 9);
  assign w578[44] = |(datain[135:132] ^ 0);
  assign w578[45] = |(datain[131:128] ^ 4);
  assign w578[46] = |(datain[127:124] ^ 0);
  assign w578[47] = |(datain[123:120] ^ 0);
  assign w578[48] = |(datain[119:116] ^ 15);
  assign w578[49] = |(datain[115:112] ^ 12);
  assign w578[50] = |(datain[111:108] ^ 15);
  assign w578[51] = |(datain[107:104] ^ 3);
  assign w578[52] = |(datain[103:100] ^ 10);
  assign w578[53] = |(datain[99:96] ^ 4);
  assign w578[54] = |(datain[95:92] ^ 11);
  assign w578[55] = |(datain[91:88] ^ 4);
  assign w578[56] = |(datain[87:84] ^ 1);
  assign w578[57] = |(datain[83:80] ^ 10);
  assign w578[58] = |(datain[79:76] ^ 8);
  assign w578[59] = |(datain[75:72] ^ 13);
  assign comp[578] = ~(|w578);
  wire [74-1:0] w579;
  assign w579[0] = |(datain[311:308] ^ 0);
  assign w579[1] = |(datain[307:304] ^ 4);
  assign w579[2] = |(datain[303:300] ^ 0);
  assign w579[3] = |(datain[299:296] ^ 0);
  assign w579[4] = |(datain[295:292] ^ 8);
  assign w579[5] = |(datain[291:288] ^ 13);
  assign w579[6] = |(datain[287:284] ^ 9);
  assign w579[7] = |(datain[283:280] ^ 6);
  assign w579[8] = |(datain[279:276] ^ 15);
  assign w579[9] = |(datain[275:272] ^ 11);
  assign w579[10] = |(datain[271:268] ^ 0);
  assign w579[11] = |(datain[267:264] ^ 1);
  assign w579[12] = |(datain[263:260] ^ 12);
  assign w579[13] = |(datain[259:256] ^ 13);
  assign w579[14] = |(datain[255:252] ^ 2);
  assign w579[15] = |(datain[251:248] ^ 1);
  assign w579[16] = |(datain[247:244] ^ 11);
  assign w579[17] = |(datain[243:240] ^ 8);
  assign w579[18] = |(datain[239:236] ^ 0);
  assign w579[19] = |(datain[235:232] ^ 2);
  assign w579[20] = |(datain[231:228] ^ 4);
  assign w579[21] = |(datain[227:224] ^ 2);
  assign w579[22] = |(datain[223:220] ^ 3);
  assign w579[23] = |(datain[219:216] ^ 3);
  assign w579[24] = |(datain[215:212] ^ 12);
  assign w579[25] = |(datain[211:208] ^ 9);
  assign w579[26] = |(datain[207:204] ^ 3);
  assign w579[27] = |(datain[203:200] ^ 3);
  assign w579[28] = |(datain[199:196] ^ 13);
  assign w579[29] = |(datain[195:192] ^ 2);
  assign w579[30] = |(datain[191:188] ^ 12);
  assign w579[31] = |(datain[187:184] ^ 13);
  assign w579[32] = |(datain[183:180] ^ 2);
  assign w579[33] = |(datain[179:176] ^ 1);
  assign w579[34] = |(datain[175:172] ^ 11);
  assign w579[35] = |(datain[171:168] ^ 4);
  assign w579[36] = |(datain[167:164] ^ 4);
  assign w579[37] = |(datain[163:160] ^ 0);
  assign w579[38] = |(datain[159:156] ^ 8);
  assign w579[39] = |(datain[155:152] ^ 11);
  assign w579[40] = |(datain[151:148] ^ 0);
  assign w579[41] = |(datain[147:144] ^ 14);
  assign w579[42] = |(datain[143:140] ^ 3);
  assign w579[43] = |(datain[139:136] ^ 12);
  assign w579[44] = |(datain[135:132] ^ 0);
  assign w579[45] = |(datain[131:128] ^ 2);
  assign w579[46] = |(datain[127:124] ^ 11);
  assign w579[47] = |(datain[123:120] ^ 10);
  assign w579[48] = |(datain[119:116] ^ 0);
  assign w579[49] = |(datain[115:112] ^ 4);
  assign w579[50] = |(datain[111:108] ^ 0);
  assign w579[51] = |(datain[107:104] ^ 1);
  assign w579[52] = |(datain[103:100] ^ 12);
  assign w579[53] = |(datain[99:96] ^ 13);
  assign w579[54] = |(datain[95:92] ^ 2);
  assign w579[55] = |(datain[91:88] ^ 1);
  assign w579[56] = |(datain[87:84] ^ 11);
  assign w579[57] = |(datain[83:80] ^ 8);
  assign w579[58] = |(datain[79:76] ^ 0);
  assign w579[59] = |(datain[75:72] ^ 1);
  assign w579[60] = |(datain[71:68] ^ 4);
  assign w579[61] = |(datain[67:64] ^ 3);
  assign w579[62] = |(datain[63:60] ^ 8);
  assign w579[63] = |(datain[59:56] ^ 11);
  assign w579[64] = |(datain[55:52] ^ 8);
  assign w579[65] = |(datain[51:48] ^ 14);
  assign w579[66] = |(datain[47:44] ^ 2);
  assign w579[67] = |(datain[43:40] ^ 15);
  assign w579[68] = |(datain[39:36] ^ 0);
  assign w579[69] = |(datain[35:32] ^ 2);
  assign w579[70] = |(datain[31:28] ^ 12);
  assign w579[71] = |(datain[27:24] ^ 13);
  assign w579[72] = |(datain[23:20] ^ 2);
  assign w579[73] = |(datain[19:16] ^ 1);
  assign comp[579] = ~(|w579);
  wire [74-1:0] w580;
  assign w580[0] = |(datain[311:308] ^ 1);
  assign w580[1] = |(datain[307:304] ^ 15);
  assign w580[2] = |(datain[303:300] ^ 0);
  assign w580[3] = |(datain[299:296] ^ 2);
  assign w580[4] = |(datain[295:292] ^ 12);
  assign w580[5] = |(datain[291:288] ^ 6);
  assign w580[6] = |(datain[287:284] ^ 8);
  assign w580[7] = |(datain[283:280] ^ 6);
  assign w580[8] = |(datain[279:276] ^ 2);
  assign w580[9] = |(datain[275:272] ^ 0);
  assign w580[10] = |(datain[271:268] ^ 0);
  assign w580[11] = |(datain[267:264] ^ 2);
  assign w580[12] = |(datain[263:260] ^ 13);
  assign w580[13] = |(datain[259:256] ^ 14);
  assign w580[14] = |(datain[255:252] ^ 11);
  assign w580[15] = |(datain[251:248] ^ 4);
  assign w580[16] = |(datain[247:244] ^ 4);
  assign w580[17] = |(datain[243:240] ^ 2);
  assign w580[18] = |(datain[239:236] ^ 11);
  assign w580[19] = |(datain[235:232] ^ 0);
  assign w580[20] = |(datain[231:228] ^ 0);
  assign w580[21] = |(datain[227:224] ^ 0);
  assign w580[22] = |(datain[223:220] ^ 3);
  assign w580[23] = |(datain[219:216] ^ 3);
  assign w580[24] = |(datain[215:212] ^ 12);
  assign w580[25] = |(datain[211:208] ^ 9);
  assign w580[26] = |(datain[207:204] ^ 3);
  assign w580[27] = |(datain[203:200] ^ 3);
  assign w580[28] = |(datain[199:196] ^ 13);
  assign w580[29] = |(datain[195:192] ^ 2);
  assign w580[30] = |(datain[191:188] ^ 12);
  assign w580[31] = |(datain[187:184] ^ 13);
  assign w580[32] = |(datain[183:180] ^ 2);
  assign w580[33] = |(datain[179:176] ^ 1);
  assign w580[34] = |(datain[175:172] ^ 11);
  assign w580[35] = |(datain[171:168] ^ 4);
  assign w580[36] = |(datain[167:164] ^ 4);
  assign w580[37] = |(datain[163:160] ^ 0);
  assign w580[38] = |(datain[159:156] ^ 11);
  assign w580[39] = |(datain[155:152] ^ 9);
  assign w580[40] = |(datain[151:148] ^ 0);
  assign w580[41] = |(datain[147:144] ^ 4);
  assign w580[42] = |(datain[143:140] ^ 0);
  assign w580[43] = |(datain[139:136] ^ 0);
  assign w580[44] = |(datain[135:132] ^ 8);
  assign w580[45] = |(datain[131:128] ^ 13);
  assign w580[46] = |(datain[127:124] ^ 9);
  assign w580[47] = |(datain[123:120] ^ 6);
  assign w580[48] = |(datain[119:116] ^ 1);
  assign w580[49] = |(datain[115:112] ^ 13);
  assign w580[50] = |(datain[111:108] ^ 0);
  assign w580[51] = |(datain[107:104] ^ 2);
  assign w580[52] = |(datain[103:100] ^ 12);
  assign w580[53] = |(datain[99:96] ^ 13);
  assign w580[54] = |(datain[95:92] ^ 2);
  assign w580[55] = |(datain[91:88] ^ 1);
  assign w580[56] = |(datain[87:84] ^ 11);
  assign w580[57] = |(datain[83:80] ^ 4);
  assign w580[58] = |(datain[79:76] ^ 4);
  assign w580[59] = |(datain[75:72] ^ 2);
  assign w580[60] = |(datain[71:68] ^ 11);
  assign w580[61] = |(datain[67:64] ^ 0);
  assign w580[62] = |(datain[63:60] ^ 0);
  assign w580[63] = |(datain[59:56] ^ 2);
  assign w580[64] = |(datain[55:52] ^ 3);
  assign w580[65] = |(datain[51:48] ^ 3);
  assign w580[66] = |(datain[47:44] ^ 12);
  assign w580[67] = |(datain[43:40] ^ 9);
  assign w580[68] = |(datain[39:36] ^ 3);
  assign w580[69] = |(datain[35:32] ^ 3);
  assign w580[70] = |(datain[31:28] ^ 13);
  assign w580[71] = |(datain[27:24] ^ 2);
  assign w580[72] = |(datain[23:20] ^ 12);
  assign w580[73] = |(datain[19:16] ^ 13);
  assign comp[580] = ~(|w580);
  wire [42-1:0] w581;
  assign w581[0] = |(datain[311:308] ^ 0);
  assign w581[1] = |(datain[307:304] ^ 1);
  assign w581[2] = |(datain[303:300] ^ 11);
  assign w581[3] = |(datain[299:296] ^ 15);
  assign w581[4] = |(datain[295:292] ^ 0);
  assign w581[5] = |(datain[291:288] ^ 0);
  assign w581[6] = |(datain[287:284] ^ 0);
  assign w581[7] = |(datain[283:280] ^ 1);
  assign w581[8] = |(datain[279:276] ^ 11);
  assign w581[9] = |(datain[275:272] ^ 9);
  assign w581[10] = |(datain[271:268] ^ 0);
  assign w581[11] = |(datain[267:264] ^ 4);
  assign w581[12] = |(datain[263:260] ^ 0);
  assign w581[13] = |(datain[259:256] ^ 0);
  assign w581[14] = |(datain[255:252] ^ 15);
  assign w581[15] = |(datain[251:248] ^ 12);
  assign w581[16] = |(datain[247:244] ^ 15);
  assign w581[17] = |(datain[243:240] ^ 3);
  assign w581[18] = |(datain[239:236] ^ 10);
  assign w581[19] = |(datain[235:232] ^ 4);
  assign w581[20] = |(datain[231:228] ^ 11);
  assign w581[21] = |(datain[227:224] ^ 4);
  assign w581[22] = |(datain[223:220] ^ 1);
  assign w581[23] = |(datain[219:216] ^ 10);
  assign w581[24] = |(datain[215:212] ^ 8);
  assign w581[25] = |(datain[211:208] ^ 13);
  assign w581[26] = |(datain[207:204] ^ 9);
  assign w581[27] = |(datain[203:200] ^ 6);
  assign w581[28] = |(datain[199:196] ^ 11);
  assign w581[29] = |(datain[195:192] ^ 14);
  assign w581[30] = |(datain[191:188] ^ 0);
  assign w581[31] = |(datain[187:184] ^ 2);
  assign w581[32] = |(datain[183:180] ^ 12);
  assign w581[33] = |(datain[179:176] ^ 13);
  assign w581[34] = |(datain[175:172] ^ 2);
  assign w581[35] = |(datain[171:168] ^ 1);
  assign w581[36] = |(datain[167:164] ^ 11);
  assign w581[37] = |(datain[163:160] ^ 4);
  assign w581[38] = |(datain[159:156] ^ 4);
  assign w581[39] = |(datain[155:152] ^ 14);
  assign w581[40] = |(datain[151:148] ^ 8);
  assign w581[41] = |(datain[147:144] ^ 13);
  assign comp[581] = ~(|w581);
  wire [42-1:0] w582;
  assign w582[0] = |(datain[311:308] ^ 0);
  assign w582[1] = |(datain[307:304] ^ 1);
  assign w582[2] = |(datain[303:300] ^ 11);
  assign w582[3] = |(datain[299:296] ^ 15);
  assign w582[4] = |(datain[295:292] ^ 0);
  assign w582[5] = |(datain[291:288] ^ 0);
  assign w582[6] = |(datain[287:284] ^ 0);
  assign w582[7] = |(datain[283:280] ^ 1);
  assign w582[8] = |(datain[279:276] ^ 11);
  assign w582[9] = |(datain[275:272] ^ 9);
  assign w582[10] = |(datain[271:268] ^ 0);
  assign w582[11] = |(datain[267:264] ^ 4);
  assign w582[12] = |(datain[263:260] ^ 0);
  assign w582[13] = |(datain[259:256] ^ 0);
  assign w582[14] = |(datain[255:252] ^ 15);
  assign w582[15] = |(datain[251:248] ^ 12);
  assign w582[16] = |(datain[247:244] ^ 15);
  assign w582[17] = |(datain[243:240] ^ 3);
  assign w582[18] = |(datain[239:236] ^ 10);
  assign w582[19] = |(datain[235:232] ^ 4);
  assign w582[20] = |(datain[231:228] ^ 11);
  assign w582[21] = |(datain[227:224] ^ 4);
  assign w582[22] = |(datain[223:220] ^ 1);
  assign w582[23] = |(datain[219:216] ^ 10);
  assign w582[24] = |(datain[215:212] ^ 8);
  assign w582[25] = |(datain[211:208] ^ 13);
  assign w582[26] = |(datain[207:204] ^ 9);
  assign w582[27] = |(datain[203:200] ^ 6);
  assign w582[28] = |(datain[199:196] ^ 12);
  assign w582[29] = |(datain[195:192] ^ 6);
  assign w582[30] = |(datain[191:188] ^ 0);
  assign w582[31] = |(datain[187:184] ^ 2);
  assign w582[32] = |(datain[183:180] ^ 12);
  assign w582[33] = |(datain[179:176] ^ 13);
  assign w582[34] = |(datain[175:172] ^ 2);
  assign w582[35] = |(datain[171:168] ^ 1);
  assign w582[36] = |(datain[167:164] ^ 11);
  assign w582[37] = |(datain[163:160] ^ 4);
  assign w582[38] = |(datain[159:156] ^ 4);
  assign w582[39] = |(datain[155:152] ^ 14);
  assign w582[40] = |(datain[151:148] ^ 8);
  assign w582[41] = |(datain[147:144] ^ 13);
  assign comp[582] = ~(|w582);
  wire [46-1:0] w583;
  assign w583[0] = |(datain[311:308] ^ 11);
  assign w583[1] = |(datain[307:304] ^ 6);
  assign w583[2] = |(datain[303:300] ^ 0);
  assign w583[3] = |(datain[299:296] ^ 5);
  assign w583[4] = |(datain[295:292] ^ 0);
  assign w583[5] = |(datain[291:288] ^ 1);
  assign w583[6] = |(datain[287:284] ^ 11);
  assign w583[7] = |(datain[283:280] ^ 15);
  assign w583[8] = |(datain[279:276] ^ 0);
  assign w583[9] = |(datain[275:272] ^ 0);
  assign w583[10] = |(datain[271:268] ^ 0);
  assign w583[11] = |(datain[267:264] ^ 1);
  assign w583[12] = |(datain[263:260] ^ 11);
  assign w583[13] = |(datain[259:256] ^ 9);
  assign w583[14] = |(datain[255:252] ^ 0);
  assign w583[15] = |(datain[251:248] ^ 4);
  assign w583[16] = |(datain[247:244] ^ 0);
  assign w583[17] = |(datain[243:240] ^ 0);
  assign w583[18] = |(datain[239:236] ^ 15);
  assign w583[19] = |(datain[235:232] ^ 12);
  assign w583[20] = |(datain[231:228] ^ 15);
  assign w583[21] = |(datain[227:224] ^ 3);
  assign w583[22] = |(datain[223:220] ^ 10);
  assign w583[23] = |(datain[219:216] ^ 4);
  assign w583[24] = |(datain[215:212] ^ 11);
  assign w583[25] = |(datain[211:208] ^ 4);
  assign w583[26] = |(datain[207:204] ^ 1);
  assign w583[27] = |(datain[203:200] ^ 10);
  assign w583[28] = |(datain[199:196] ^ 8);
  assign w583[29] = |(datain[195:192] ^ 13);
  assign w583[30] = |(datain[191:188] ^ 9);
  assign w583[31] = |(datain[187:184] ^ 6);
  assign w583[32] = |(datain[183:180] ^ 12);
  assign w583[33] = |(datain[179:176] ^ 8);
  assign w583[34] = |(datain[175:172] ^ 0);
  assign w583[35] = |(datain[171:168] ^ 2);
  assign w583[36] = |(datain[167:164] ^ 12);
  assign w583[37] = |(datain[163:160] ^ 13);
  assign w583[38] = |(datain[159:156] ^ 2);
  assign w583[39] = |(datain[155:152] ^ 1);
  assign w583[40] = |(datain[151:148] ^ 11);
  assign w583[41] = |(datain[147:144] ^ 4);
  assign w583[42] = |(datain[143:140] ^ 4);
  assign w583[43] = |(datain[139:136] ^ 14);
  assign w583[44] = |(datain[135:132] ^ 8);
  assign w583[45] = |(datain[131:128] ^ 13);
  assign comp[583] = ~(|w583);
  wire [42-1:0] w584;
  assign w584[0] = |(datain[311:308] ^ 5);
  assign w584[1] = |(datain[307:304] ^ 13);
  assign w584[2] = |(datain[303:300] ^ 8);
  assign w584[3] = |(datain[299:296] ^ 1);
  assign w584[4] = |(datain[295:292] ^ 14);
  assign w584[5] = |(datain[291:288] ^ 13);
  assign w584[6] = |(datain[287:284] ^ 0);
  assign w584[7] = |(datain[283:280] ^ 11);
  assign w584[8] = |(datain[279:276] ^ 0);
  assign w584[9] = |(datain[275:272] ^ 1);
  assign w584[10] = |(datain[271:268] ^ 8);
  assign w584[11] = |(datain[267:264] ^ 13);
  assign w584[12] = |(datain[263:260] ^ 9);
  assign w584[13] = |(datain[259:256] ^ 14);
  assign w584[14] = |(datain[255:252] ^ 2);
  assign w584[15] = |(datain[251:248] ^ 10);
  assign w584[16] = |(datain[247:244] ^ 0);
  assign w584[17] = |(datain[243:240] ^ 1);
  assign w584[18] = |(datain[239:236] ^ 5);
  assign w584[19] = |(datain[235:232] ^ 3);
  assign w584[20] = |(datain[231:228] ^ 8);
  assign w584[21] = |(datain[227:224] ^ 10);
  assign w584[22] = |(datain[223:220] ^ 8);
  assign w584[23] = |(datain[219:216] ^ 6);
  assign w584[24] = |(datain[215:212] ^ 2);
  assign w584[25] = |(datain[211:208] ^ 2);
  assign w584[26] = |(datain[207:204] ^ 0);
  assign w584[27] = |(datain[203:200] ^ 1);
  assign w584[28] = |(datain[199:196] ^ 11);
  assign w584[29] = |(datain[195:192] ^ 9);
  assign w584[30] = |(datain[191:188] ^ 10);
  assign w584[31] = |(datain[187:184] ^ 2);
  assign w584[32] = |(datain[183:180] ^ 0);
  assign w584[33] = |(datain[179:176] ^ 2);
  assign w584[34] = |(datain[175:172] ^ 3);
  assign w584[35] = |(datain[171:168] ^ 0);
  assign w584[36] = |(datain[167:164] ^ 0);
  assign w584[37] = |(datain[163:160] ^ 7);
  assign w584[38] = |(datain[159:156] ^ 4);
  assign w584[39] = |(datain[155:152] ^ 3);
  assign w584[40] = |(datain[151:148] ^ 14);
  assign w584[41] = |(datain[147:144] ^ 2);
  assign comp[584] = ~(|w584);
  wire [48-1:0] w585;
  assign w585[0] = |(datain[311:308] ^ 14);
  assign w585[1] = |(datain[307:304] ^ 8);
  assign w585[2] = |(datain[303:300] ^ 0);
  assign w585[3] = |(datain[299:296] ^ 0);
  assign w585[4] = |(datain[295:292] ^ 0);
  assign w585[5] = |(datain[291:288] ^ 0);
  assign w585[6] = |(datain[287:284] ^ 5);
  assign w585[7] = |(datain[283:280] ^ 13);
  assign w585[8] = |(datain[279:276] ^ 8);
  assign w585[9] = |(datain[275:272] ^ 1);
  assign w585[10] = |(datain[271:268] ^ 14);
  assign w585[11] = |(datain[267:264] ^ 13);
  assign w585[12] = |(datain[263:260] ^ 0);
  assign w585[13] = |(datain[259:256] ^ 11);
  assign w585[14] = |(datain[255:252] ^ 0);
  assign w585[15] = |(datain[251:248] ^ 1);
  assign w585[16] = |(datain[247:244] ^ 8);
  assign w585[17] = |(datain[243:240] ^ 13);
  assign w585[18] = |(datain[239:236] ^ 9);
  assign w585[19] = |(datain[235:232] ^ 14);
  assign w585[20] = |(datain[231:228] ^ 2);
  assign w585[21] = |(datain[227:224] ^ 11);
  assign w585[22] = |(datain[223:220] ^ 0);
  assign w585[23] = |(datain[219:216] ^ 1);
  assign w585[24] = |(datain[215:212] ^ 5);
  assign w585[25] = |(datain[211:208] ^ 3);
  assign w585[26] = |(datain[207:204] ^ 3);
  assign w585[27] = |(datain[203:200] ^ 14);
  assign w585[28] = |(datain[199:196] ^ 8);
  assign w585[29] = |(datain[195:192] ^ 10);
  assign w585[30] = |(datain[191:188] ^ 8);
  assign w585[31] = |(datain[187:184] ^ 6);
  assign w585[32] = |(datain[183:180] ^ 2);
  assign w585[33] = |(datain[179:176] ^ 3);
  assign w585[34] = |(datain[175:172] ^ 0);
  assign w585[35] = |(datain[171:168] ^ 1);
  assign w585[36] = |(datain[167:164] ^ 11);
  assign w585[37] = |(datain[163:160] ^ 9);
  assign w585[38] = |(datain[159:156] ^ 11);
  assign w585[39] = |(datain[155:152] ^ 10);
  assign w585[40] = |(datain[151:148] ^ 0);
  assign w585[41] = |(datain[147:144] ^ 2);
  assign w585[42] = |(datain[143:140] ^ 3);
  assign w585[43] = |(datain[139:136] ^ 0);
  assign w585[44] = |(datain[135:132] ^ 0);
  assign w585[45] = |(datain[131:128] ^ 7);
  assign w585[46] = |(datain[127:124] ^ 4);
  assign w585[47] = |(datain[123:120] ^ 3);
  assign comp[585] = ~(|w585);
  wire [42-1:0] w586;
  assign w586[0] = |(datain[311:308] ^ 0);
  assign w586[1] = |(datain[307:304] ^ 1);
  assign w586[2] = |(datain[303:300] ^ 11);
  assign w586[3] = |(datain[299:296] ^ 15);
  assign w586[4] = |(datain[295:292] ^ 0);
  assign w586[5] = |(datain[291:288] ^ 0);
  assign w586[6] = |(datain[287:284] ^ 0);
  assign w586[7] = |(datain[283:280] ^ 1);
  assign w586[8] = |(datain[279:276] ^ 11);
  assign w586[9] = |(datain[275:272] ^ 9);
  assign w586[10] = |(datain[271:268] ^ 0);
  assign w586[11] = |(datain[267:264] ^ 4);
  assign w586[12] = |(datain[263:260] ^ 0);
  assign w586[13] = |(datain[259:256] ^ 0);
  assign w586[14] = |(datain[255:252] ^ 15);
  assign w586[15] = |(datain[251:248] ^ 12);
  assign w586[16] = |(datain[247:244] ^ 15);
  assign w586[17] = |(datain[243:240] ^ 3);
  assign w586[18] = |(datain[239:236] ^ 10);
  assign w586[19] = |(datain[235:232] ^ 4);
  assign w586[20] = |(datain[231:228] ^ 11);
  assign w586[21] = |(datain[227:224] ^ 4);
  assign w586[22] = |(datain[223:220] ^ 1);
  assign w586[23] = |(datain[219:216] ^ 10);
  assign w586[24] = |(datain[215:212] ^ 8);
  assign w586[25] = |(datain[211:208] ^ 13);
  assign w586[26] = |(datain[207:204] ^ 9);
  assign w586[27] = |(datain[203:200] ^ 6);
  assign w586[28] = |(datain[199:196] ^ 14);
  assign w586[29] = |(datain[195:192] ^ 11);
  assign w586[30] = |(datain[191:188] ^ 0);
  assign w586[31] = |(datain[187:184] ^ 3);
  assign w586[32] = |(datain[183:180] ^ 12);
  assign w586[33] = |(datain[179:176] ^ 13);
  assign w586[34] = |(datain[175:172] ^ 2);
  assign w586[35] = |(datain[171:168] ^ 1);
  assign w586[36] = |(datain[167:164] ^ 11);
  assign w586[37] = |(datain[163:160] ^ 4);
  assign w586[38] = |(datain[159:156] ^ 4);
  assign w586[39] = |(datain[155:152] ^ 14);
  assign w586[40] = |(datain[151:148] ^ 8);
  assign w586[41] = |(datain[147:144] ^ 13);
  assign comp[586] = ~(|w586);
  wire [44-1:0] w587;
  assign w587[0] = |(datain[311:308] ^ 11);
  assign w587[1] = |(datain[307:304] ^ 9);
  assign w587[2] = |(datain[303:300] ^ 0);
  assign w587[3] = |(datain[299:296] ^ 4);
  assign w587[4] = |(datain[295:292] ^ 0);
  assign w587[5] = |(datain[291:288] ^ 0);
  assign w587[6] = |(datain[287:284] ^ 8);
  assign w587[7] = |(datain[283:280] ^ 13);
  assign w587[8] = |(datain[279:276] ^ 9);
  assign w587[9] = |(datain[275:272] ^ 6);
  assign w587[10] = |(datain[271:268] ^ 0);
  assign w587[11] = |(datain[267:264] ^ 4);
  assign w587[12] = |(datain[263:260] ^ 0);
  assign w587[13] = |(datain[259:256] ^ 1);
  assign w587[14] = |(datain[255:252] ^ 12);
  assign w587[15] = |(datain[251:248] ^ 13);
  assign w587[16] = |(datain[247:244] ^ 2);
  assign w587[17] = |(datain[243:240] ^ 1);
  assign w587[18] = |(datain[239:236] ^ 8);
  assign w587[19] = |(datain[235:232] ^ 0);
  assign w587[20] = |(datain[231:228] ^ 11);
  assign w587[21] = |(datain[227:224] ^ 14);
  assign w587[22] = |(datain[223:220] ^ 0);
  assign w587[23] = |(datain[219:216] ^ 7);
  assign w587[24] = |(datain[215:212] ^ 0);
  assign w587[25] = |(datain[211:208] ^ 1);
  assign w587[26] = |(datain[207:204] ^ 1);
  assign w587[27] = |(datain[203:200] ^ 10);
  assign w587[28] = |(datain[199:196] ^ 7);
  assign w587[29] = |(datain[195:192] ^ 4);
  assign w587[30] = |(datain[191:188] ^ 12);
  assign w587[31] = |(datain[187:184] ^ 10);
  assign w587[32] = |(datain[183:180] ^ 8);
  assign w587[33] = |(datain[179:176] ^ 0);
  assign w587[34] = |(datain[175:172] ^ 11);
  assign w587[35] = |(datain[171:168] ^ 14);
  assign w587[36] = |(datain[167:164] ^ 0);
  assign w587[37] = |(datain[163:160] ^ 4);
  assign w587[38] = |(datain[159:156] ^ 0);
  assign w587[39] = |(datain[155:152] ^ 1);
  assign w587[40] = |(datain[151:148] ^ 4);
  assign w587[41] = |(datain[147:144] ^ 13);
  assign w587[42] = |(datain[143:140] ^ 7);
  assign w587[43] = |(datain[139:136] ^ 4);
  assign comp[587] = ~(|w587);
  wire [32-1:0] w588;
  assign w588[0] = |(datain[311:308] ^ 4);
  assign w588[1] = |(datain[307:304] ^ 13);
  assign w588[2] = |(datain[303:300] ^ 0);
  assign w588[3] = |(datain[299:296] ^ 0);
  assign w588[4] = |(datain[295:292] ^ 8);
  assign w588[5] = |(datain[291:288] ^ 1);
  assign w588[6] = |(datain[287:284] ^ 12);
  assign w588[7] = |(datain[283:280] ^ 3);
  assign w588[8] = |(datain[279:276] ^ 0);
  assign w588[9] = |(datain[275:272] ^ 0);
  assign w588[10] = |(datain[271:268] ^ 0);
  assign w588[11] = |(datain[267:264] ^ 2);
  assign w588[12] = |(datain[263:260] ^ 14);
  assign w588[13] = |(datain[259:256] ^ 2);
  assign w588[14] = |(datain[255:252] ^ 15);
  assign w588[15] = |(datain[251:248] ^ 4);
  assign w588[16] = |(datain[247:244] ^ 10);
  assign w588[17] = |(datain[243:240] ^ 1);
  assign w588[18] = |(datain[239:236] ^ 1);
  assign w588[19] = |(datain[235:232] ^ 3);
  assign w588[20] = |(datain[231:228] ^ 0);
  assign w588[21] = |(datain[227:224] ^ 4);
  assign w588[22] = |(datain[223:220] ^ 2);
  assign w588[23] = |(datain[219:216] ^ 13);
  assign w588[24] = |(datain[215:212] ^ 0);
  assign w588[25] = |(datain[211:208] ^ 7);
  assign w588[26] = |(datain[207:204] ^ 0);
  assign w588[27] = |(datain[203:200] ^ 0);
  assign w588[28] = |(datain[199:196] ^ 10);
  assign w588[29] = |(datain[195:192] ^ 3);
  assign w588[30] = |(datain[191:188] ^ 1);
  assign w588[31] = |(datain[187:184] ^ 3);
  assign comp[588] = ~(|w588);
  wire [32-1:0] w589;
  assign w589[0] = |(datain[311:308] ^ 10);
  assign w589[1] = |(datain[307:304] ^ 0);
  assign w589[2] = |(datain[303:300] ^ 0);
  assign w589[3] = |(datain[299:296] ^ 6);
  assign w589[4] = |(datain[295:292] ^ 7);
  assign w589[5] = |(datain[291:288] ^ 12);
  assign w589[6] = |(datain[287:284] ^ 10);
  assign w589[7] = |(datain[283:280] ^ 2);
  assign w589[8] = |(datain[279:276] ^ 0);
  assign w589[9] = |(datain[275:272] ^ 9);
  assign w589[10] = |(datain[271:268] ^ 7);
  assign w589[11] = |(datain[267:264] ^ 12);
  assign w589[12] = |(datain[263:260] ^ 8);
  assign w589[13] = |(datain[259:256] ^ 11);
  assign w589[14] = |(datain[255:252] ^ 0);
  assign w589[15] = |(datain[251:248] ^ 14);
  assign w589[16] = |(datain[247:244] ^ 0);
  assign w589[17] = |(datain[243:240] ^ 7);
  assign w589[18] = |(datain[239:236] ^ 7);
  assign w589[19] = |(datain[235:232] ^ 12);
  assign w589[20] = |(datain[231:228] ^ 8);
  assign w589[21] = |(datain[227:224] ^ 9);
  assign w589[22] = |(datain[223:220] ^ 0);
  assign w589[23] = |(datain[219:216] ^ 14);
  assign w589[24] = |(datain[215:212] ^ 0);
  assign w589[25] = |(datain[211:208] ^ 10);
  assign w589[26] = |(datain[207:204] ^ 7);
  assign w589[27] = |(datain[203:200] ^ 12);
  assign w589[28] = |(datain[199:196] ^ 14);
  assign w589[29] = |(datain[195:192] ^ 8);
  assign w589[30] = |(datain[191:188] ^ 5);
  assign w589[31] = |(datain[187:184] ^ 9);
  assign comp[589] = ~(|w589);
  wire [52-1:0] w590;
  assign w590[0] = |(datain[311:308] ^ 14);
  assign w590[1] = |(datain[307:304] ^ 8);
  assign w590[2] = |(datain[303:300] ^ 0);
  assign w590[3] = |(datain[299:296] ^ 0);
  assign w590[4] = |(datain[295:292] ^ 0);
  assign w590[5] = |(datain[291:288] ^ 0);
  assign w590[6] = |(datain[287:284] ^ 5);
  assign w590[7] = |(datain[283:280] ^ 11);
  assign w590[8] = |(datain[279:276] ^ 5);
  assign w590[9] = |(datain[275:272] ^ 3);
  assign w590[10] = |(datain[271:268] ^ 8);
  assign w590[11] = |(datain[267:264] ^ 3);
  assign w590[12] = |(datain[263:260] ^ 12);
  assign w590[13] = |(datain[259:256] ^ 3);
  assign w590[14] = |(datain[255:252] ^ 1);
  assign w590[15] = |(datain[251:248] ^ 7);
  assign w590[16] = |(datain[247:244] ^ 9);
  assign w590[17] = |(datain[243:240] ^ 0);
  assign w590[18] = |(datain[239:236] ^ 11);
  assign w590[19] = |(datain[235:232] ^ 10);
  assign w590[20] = |(datain[231:228] ^ 0);
  assign w590[21] = |(datain[227:224] ^ 0);
  assign w590[22] = |(datain[223:220] ^ 0);
  assign w590[23] = |(datain[219:216] ^ 0);
  assign w590[24] = |(datain[215:212] ^ 11);
  assign w590[25] = |(datain[211:208] ^ 9);
  assign w590[26] = |(datain[207:204] ^ 15);
  assign w590[27] = |(datain[203:200] ^ 4);
  assign w590[28] = |(datain[199:196] ^ 0);
  assign w590[29] = |(datain[195:192] ^ 1);
  assign w590[30] = |(datain[191:188] ^ 2);
  assign w590[31] = |(datain[187:184] ^ 14);
  assign w590[32] = |(datain[183:180] ^ 3);
  assign w590[33] = |(datain[179:176] ^ 1);
  assign w590[34] = |(datain[175:172] ^ 1);
  assign w590[35] = |(datain[171:168] ^ 7);
  assign w590[36] = |(datain[167:164] ^ 14);
  assign w590[37] = |(datain[163:160] ^ 3);
  assign w590[38] = |(datain[159:156] ^ 0);
  assign w590[39] = |(datain[155:152] ^ 6);
  assign w590[40] = |(datain[151:148] ^ 4);
  assign w590[41] = |(datain[147:144] ^ 3);
  assign w590[42] = |(datain[143:140] ^ 4);
  assign w590[43] = |(datain[139:136] ^ 3);
  assign w590[44] = |(datain[135:132] ^ 4);
  assign w590[45] = |(datain[131:128] ^ 9);
  assign w590[46] = |(datain[127:124] ^ 4);
  assign w590[47] = |(datain[123:120] ^ 9);
  assign w590[48] = |(datain[119:116] ^ 14);
  assign w590[49] = |(datain[115:112] ^ 11);
  assign w590[50] = |(datain[111:108] ^ 15);
  assign w590[51] = |(datain[107:104] ^ 5);
  assign comp[590] = ~(|w590);
  wire [76-1:0] w591;
  assign w591[0] = |(datain[311:308] ^ 0);
  assign w591[1] = |(datain[307:304] ^ 14);
  assign w591[2] = |(datain[303:300] ^ 1);
  assign w591[3] = |(datain[299:296] ^ 3);
  assign w591[4] = |(datain[295:292] ^ 0);
  assign w591[5] = |(datain[291:288] ^ 4);
  assign w591[6] = |(datain[287:284] ^ 10);
  assign w591[7] = |(datain[283:280] ^ 1);
  assign w591[8] = |(datain[279:276] ^ 1);
  assign w591[9] = |(datain[275:272] ^ 3);
  assign w591[10] = |(datain[271:268] ^ 0);
  assign w591[11] = |(datain[267:264] ^ 4);
  assign w591[12] = |(datain[263:260] ^ 12);
  assign w591[13] = |(datain[259:256] ^ 1);
  assign w591[14] = |(datain[255:252] ^ 14);
  assign w591[15] = |(datain[251:248] ^ 0);
  assign w591[16] = |(datain[247:244] ^ 0);
  assign w591[17] = |(datain[243:240] ^ 6);
  assign w591[18] = |(datain[239:236] ^ 8);
  assign w591[19] = |(datain[235:232] ^ 14);
  assign w591[20] = |(datain[231:228] ^ 12);
  assign w591[21] = |(datain[227:224] ^ 0);
  assign w591[22] = |(datain[223:220] ^ 1);
  assign w591[23] = |(datain[219:216] ^ 14);
  assign w591[24] = |(datain[215:212] ^ 5);
  assign w591[25] = |(datain[211:208] ^ 6);
  assign w591[26] = |(datain[207:204] ^ 0);
  assign w591[27] = |(datain[203:200] ^ 6);
  assign w591[28] = |(datain[199:196] ^ 6);
  assign w591[29] = |(datain[195:192] ^ 8);
  assign w591[30] = |(datain[191:188] ^ 3);
  assign w591[31] = |(datain[187:184] ^ 8);
  assign w591[32] = |(datain[183:180] ^ 0);
  assign w591[33] = |(datain[179:176] ^ 0);
  assign w591[34] = |(datain[175:172] ^ 3);
  assign w591[35] = |(datain[171:168] ^ 3);
  assign w591[36] = |(datain[167:164] ^ 15);
  assign w591[37] = |(datain[163:160] ^ 15);
  assign w591[38] = |(datain[159:156] ^ 8);
  assign w591[39] = |(datain[155:152] ^ 9);
  assign w591[40] = |(datain[151:148] ^ 12);
  assign w591[41] = |(datain[147:144] ^ 1);
  assign w591[42] = |(datain[143:140] ^ 15);
  assign w591[43] = |(datain[139:136] ^ 3);
  assign w591[44] = |(datain[135:132] ^ 10);
  assign w591[45] = |(datain[131:128] ^ 4);
  assign w591[46] = |(datain[127:124] ^ 12);
  assign w591[47] = |(datain[123:120] ^ 11);
  assign w591[48] = |(datain[119:116] ^ 12);
  assign w591[49] = |(datain[115:112] ^ 4);
  assign w591[50] = |(datain[111:108] ^ 0);
  assign w591[51] = |(datain[107:104] ^ 6);
  assign w591[52] = |(datain[103:100] ^ 4);
  assign w591[53] = |(datain[99:96] ^ 12);
  assign w591[54] = |(datain[95:92] ^ 0);
  assign w591[55] = |(datain[91:88] ^ 0);
  assign w591[56] = |(datain[87:84] ^ 2);
  assign w591[57] = |(datain[83:80] ^ 14);
  assign w591[58] = |(datain[79:76] ^ 10);
  assign w591[59] = |(datain[75:72] ^ 3);
  assign w591[60] = |(datain[71:68] ^ 7);
  assign w591[61] = |(datain[67:64] ^ 14);
  assign w591[62] = |(datain[63:60] ^ 0);
  assign w591[63] = |(datain[59:56] ^ 0);
  assign w591[64] = |(datain[55:52] ^ 2);
  assign w591[65] = |(datain[51:48] ^ 14);
  assign w591[66] = |(datain[47:44] ^ 8);
  assign w591[67] = |(datain[43:40] ^ 12);
  assign w591[68] = |(datain[39:36] ^ 0);
  assign w591[69] = |(datain[35:32] ^ 6);
  assign w591[70] = |(datain[31:28] ^ 8);
  assign w591[71] = |(datain[27:24] ^ 0);
  assign w591[72] = |(datain[23:20] ^ 0);
  assign w591[73] = |(datain[19:16] ^ 0);
  assign w591[74] = |(datain[15:12] ^ 12);
  assign w591[75] = |(datain[11:8] ^ 7);
  assign comp[591] = ~(|w591);
  wire [74-1:0] w592;
  assign w592[0] = |(datain[311:308] ^ 5);
  assign w592[1] = |(datain[307:304] ^ 8);
  assign w592[2] = |(datain[303:300] ^ 0);
  assign w592[3] = |(datain[299:296] ^ 5);
  assign w592[4] = |(datain[295:292] ^ 2);
  assign w592[5] = |(datain[291:288] ^ 7);
  assign w592[6] = |(datain[287:284] ^ 0);
  assign w592[7] = |(datain[283:280] ^ 0);
  assign w592[8] = |(datain[279:276] ^ 8);
  assign w592[9] = |(datain[275:272] ^ 11);
  assign w592[10] = |(datain[271:268] ^ 13);
  assign w592[11] = |(datain[267:264] ^ 14);
  assign w592[12] = |(datain[263:260] ^ 8);
  assign w592[13] = |(datain[259:256] ^ 1);
  assign w592[14] = |(datain[255:252] ^ 12);
  assign w592[15] = |(datain[251:248] ^ 3);
  assign w592[16] = |(datain[247:244] ^ 8);
  assign w592[17] = |(datain[243:240] ^ 6);
  assign w592[18] = |(datain[239:236] ^ 0);
  assign w592[19] = |(datain[235:232] ^ 4);
  assign w592[20] = |(datain[231:228] ^ 8);
  assign w592[21] = |(datain[227:224] ^ 11);
  assign w592[22] = |(datain[223:220] ^ 12);
  assign w592[23] = |(datain[219:216] ^ 11);
  assign w592[24] = |(datain[215:212] ^ 2);
  assign w592[25] = |(datain[211:208] ^ 11);
  assign w592[26] = |(datain[207:204] ^ 12);
  assign w592[27] = |(datain[203:200] ^ 8);
  assign w592[28] = |(datain[199:196] ^ 14);
  assign w592[29] = |(datain[195:192] ^ 8);
  assign w592[30] = |(datain[191:188] ^ 0);
  assign w592[31] = |(datain[187:184] ^ 2);
  assign w592[32] = |(datain[183:180] ^ 0);
  assign w592[33] = |(datain[179:176] ^ 0);
  assign w592[34] = |(datain[175:172] ^ 14);
  assign w592[35] = |(datain[171:168] ^ 11);
  assign w592[36] = |(datain[167:164] ^ 0);
  assign w592[37] = |(datain[163:160] ^ 11);
  assign w592[38] = |(datain[159:156] ^ 2);
  assign w592[39] = |(datain[155:152] ^ 14);
  assign w592[40] = |(datain[151:148] ^ 8);
  assign w592[41] = |(datain[147:144] ^ 10);
  assign w592[42] = |(datain[143:140] ^ 0);
  assign w592[43] = |(datain[139:136] ^ 7);
  assign w592[44] = |(datain[135:132] ^ 2);
  assign w592[45] = |(datain[131:128] ^ 14);
  assign w592[46] = |(datain[127:124] ^ 3);
  assign w592[47] = |(datain[123:120] ^ 0);
  assign w592[48] = |(datain[119:116] ^ 4);
  assign w592[49] = |(datain[115:112] ^ 7);
  assign w592[50] = |(datain[111:108] ^ 0);
  assign w592[51] = |(datain[107:104] ^ 1);
  assign w592[52] = |(datain[103:100] ^ 4);
  assign w592[53] = |(datain[99:96] ^ 11);
  assign w592[54] = |(datain[95:92] ^ 14);
  assign w592[55] = |(datain[91:88] ^ 2);
  assign w592[56] = |(datain[87:84] ^ 15);
  assign w592[57] = |(datain[83:80] ^ 6);
  assign w592[58] = |(datain[79:76] ^ 12);
  assign w592[59] = |(datain[75:72] ^ 3);
  assign w592[60] = |(datain[71:68] ^ 8);
  assign w592[61] = |(datain[67:64] ^ 3);
  assign w592[62] = |(datain[63:60] ^ 14);
  assign w592[63] = |(datain[59:56] ^ 11);
  assign w592[64] = |(datain[55:52] ^ 3);
  assign w592[65] = |(datain[51:48] ^ 6);
  assign w592[66] = |(datain[47:44] ^ 8);
  assign w592[67] = |(datain[43:40] ^ 11);
  assign w592[68] = |(datain[39:36] ^ 12);
  assign w592[69] = |(datain[35:32] ^ 11);
  assign w592[70] = |(datain[31:28] ^ 2);
  assign w592[71] = |(datain[27:24] ^ 11);
  assign w592[72] = |(datain[23:20] ^ 12);
  assign w592[73] = |(datain[19:16] ^ 14);
  assign comp[592] = ~(|w592);
  wire [74-1:0] w593;
  assign w593[0] = |(datain[311:308] ^ 5);
  assign w593[1] = |(datain[307:304] ^ 11);
  assign w593[2] = |(datain[303:300] ^ 8);
  assign w593[3] = |(datain[299:296] ^ 3);
  assign w593[4] = |(datain[295:292] ^ 12);
  assign w593[5] = |(datain[291:288] ^ 3);
  assign w593[6] = |(datain[287:284] ^ 3);
  assign w593[7] = |(datain[283:280] ^ 5);
  assign w593[8] = |(datain[279:276] ^ 8);
  assign w593[9] = |(datain[275:272] ^ 11);
  assign w593[10] = |(datain[271:268] ^ 15);
  assign w593[11] = |(datain[267:264] ^ 3);
  assign w593[12] = |(datain[263:260] ^ 8);
  assign w593[13] = |(datain[259:256] ^ 1);
  assign w593[14] = |(datain[255:252] ^ 14);
  assign w593[15] = |(datain[251:248] ^ 14);
  assign w593[16] = |(datain[247:244] ^ 7);
  assign w593[17] = |(datain[243:240] ^ 15);
  assign w593[18] = |(datain[239:236] ^ 0);
  assign w593[19] = |(datain[235:232] ^ 12);
  assign w593[20] = |(datain[231:228] ^ 15);
  assign w593[21] = |(datain[227:224] ^ 13);
  assign w593[22] = |(datain[223:220] ^ 15);
  assign w593[23] = |(datain[219:216] ^ 12);
  assign w593[24] = |(datain[215:212] ^ 0);
  assign w593[25] = |(datain[211:208] ^ 14);
  assign w593[26] = |(datain[207:204] ^ 1);
  assign w593[27] = |(datain[203:200] ^ 15);
  assign w593[28] = |(datain[199:196] ^ 11);
  assign w593[29] = |(datain[195:192] ^ 9);
  assign w593[30] = |(datain[191:188] ^ 12);
  assign w593[31] = |(datain[187:184] ^ 0);
  assign w593[32] = |(datain[183:180] ^ 0);
  assign w593[33] = |(datain[179:176] ^ 0);
  assign w593[34] = |(datain[175:172] ^ 5);
  assign w593[35] = |(datain[171:168] ^ 1);
  assign w593[36] = |(datain[167:164] ^ 11);
  assign w593[37] = |(datain[163:160] ^ 9);
  assign w593[38] = |(datain[159:156] ^ 0);
  assign w593[39] = |(datain[155:152] ^ 8);
  assign w593[40] = |(datain[151:148] ^ 0);
  assign w593[41] = |(datain[147:144] ^ 0);
  assign w593[42] = |(datain[143:140] ^ 15);
  assign w593[43] = |(datain[139:136] ^ 13);
  assign w593[44] = |(datain[135:132] ^ 15);
  assign w593[45] = |(datain[131:128] ^ 12);
  assign w593[46] = |(datain[127:124] ^ 8);
  assign w593[47] = |(datain[123:120] ^ 10);
  assign w593[48] = |(datain[119:116] ^ 1);
  assign w593[49] = |(datain[115:112] ^ 7);
  assign w593[50] = |(datain[111:108] ^ 13);
  assign w593[51] = |(datain[107:104] ^ 0);
  assign w593[52] = |(datain[103:100] ^ 13);
  assign w593[53] = |(datain[99:96] ^ 2);
  assign w593[54] = |(datain[95:92] ^ 14);
  assign w593[55] = |(datain[91:88] ^ 8);
  assign w593[56] = |(datain[87:84] ^ 0);
  assign w593[57] = |(datain[83:80] ^ 12);
  assign w593[58] = |(datain[79:76] ^ 0);
  assign w593[59] = |(datain[75:72] ^ 0);
  assign w593[60] = |(datain[71:68] ^ 4);
  assign w593[61] = |(datain[67:64] ^ 6);
  assign w593[62] = |(datain[63:60] ^ 14);
  assign w593[63] = |(datain[59:56] ^ 2);
  assign w593[64] = |(datain[55:52] ^ 15);
  assign w593[65] = |(datain[51:48] ^ 8);
  assign w593[66] = |(datain[47:44] ^ 5);
  assign w593[67] = |(datain[43:40] ^ 9);
  assign w593[68] = |(datain[39:36] ^ 4);
  assign w593[69] = |(datain[35:32] ^ 3);
  assign w593[70] = |(datain[31:28] ^ 14);
  assign w593[71] = |(datain[27:24] ^ 2);
  assign w593[72] = |(datain[23:20] ^ 14);
  assign w593[73] = |(datain[19:16] ^ 12);
  assign comp[593] = ~(|w593);
  wire [46-1:0] w594;
  assign w594[0] = |(datain[311:308] ^ 13);
  assign w594[1] = |(datain[307:304] ^ 6);
  assign w594[2] = |(datain[303:300] ^ 3);
  assign w594[3] = |(datain[299:296] ^ 1);
  assign w594[4] = |(datain[295:292] ^ 13);
  assign w594[5] = |(datain[291:288] ^ 11);
  assign w594[6] = |(datain[287:284] ^ 8);
  assign w594[7] = |(datain[283:280] ^ 14);
  assign w594[8] = |(datain[279:276] ^ 12);
  assign w594[9] = |(datain[275:272] ^ 3);
  assign w594[10] = |(datain[271:268] ^ 11);
  assign w594[11] = |(datain[267:264] ^ 11);
  assign w594[12] = |(datain[263:260] ^ 8);
  assign w594[13] = |(datain[259:256] ^ 4);
  assign w594[14] = |(datain[255:252] ^ 0);
  assign w594[15] = |(datain[251:248] ^ 0);
  assign w594[16] = |(datain[247:244] ^ 2);
  assign w594[17] = |(datain[243:240] ^ 6);
  assign w594[18] = |(datain[239:236] ^ 8);
  assign w594[19] = |(datain[235:232] ^ 11);
  assign w594[20] = |(datain[231:228] ^ 0);
  assign w594[21] = |(datain[227:224] ^ 15);
  assign w594[22] = |(datain[223:220] ^ 8);
  assign w594[23] = |(datain[219:216] ^ 9);
  assign w594[24] = |(datain[215:212] ^ 0);
  assign w594[25] = |(datain[211:208] ^ 12);
  assign w594[26] = |(datain[207:204] ^ 8);
  assign w594[27] = |(datain[203:200] ^ 9);
  assign w594[28] = |(datain[199:196] ^ 0);
  assign w594[29] = |(datain[195:192] ^ 13);
  assign w594[30] = |(datain[191:188] ^ 4);
  assign w594[31] = |(datain[187:184] ^ 6);
  assign w594[32] = |(datain[183:180] ^ 4);
  assign w594[33] = |(datain[179:176] ^ 6);
  assign w594[34] = |(datain[175:172] ^ 4);
  assign w594[35] = |(datain[171:168] ^ 7);
  assign w594[36] = |(datain[167:164] ^ 4);
  assign w594[37] = |(datain[163:160] ^ 7);
  assign w594[38] = |(datain[159:156] ^ 4);
  assign w594[39] = |(datain[155:152] ^ 3);
  assign w594[40] = |(datain[151:148] ^ 4);
  assign w594[41] = |(datain[147:144] ^ 3);
  assign w594[42] = |(datain[143:140] ^ 2);
  assign w594[43] = |(datain[139:136] ^ 6);
  assign w594[44] = |(datain[135:132] ^ 8);
  assign w594[45] = |(datain[131:128] ^ 11);
  assign comp[594] = ~(|w594);
  wire [40-1:0] w595;
  assign w595[0] = |(datain[311:308] ^ 11);
  assign w595[1] = |(datain[307:304] ^ 14);
  assign w595[2] = |(datain[303:300] ^ 0);
  assign w595[3] = |(datain[299:296] ^ 0);
  assign w595[4] = |(datain[295:292] ^ 9);
  assign w595[5] = |(datain[291:288] ^ 0);
  assign w595[6] = |(datain[287:284] ^ 8);
  assign w595[7] = |(datain[283:280] ^ 14);
  assign w595[8] = |(datain[279:276] ^ 12);
  assign w595[9] = |(datain[275:272] ^ 6);
  assign w595[10] = |(datain[271:268] ^ 2);
  assign w595[11] = |(datain[267:264] ^ 6);
  assign w595[12] = |(datain[263:260] ^ 8);
  assign w595[13] = |(datain[259:256] ^ 11);
  assign w595[14] = |(datain[255:252] ^ 0);
  assign w595[15] = |(datain[251:248] ^ 14);
  assign w595[16] = |(datain[247:244] ^ 0);
  assign w595[17] = |(datain[243:240] ^ 0);
  assign w595[18] = |(datain[239:236] ^ 9);
  assign w595[19] = |(datain[235:232] ^ 0);
  assign w595[20] = |(datain[231:228] ^ 8);
  assign w595[21] = |(datain[227:224] ^ 1);
  assign w595[22] = |(datain[223:220] ^ 15);
  assign w595[23] = |(datain[219:216] ^ 9);
  assign w595[24] = |(datain[215:212] ^ 8);
  assign w595[25] = |(datain[211:208] ^ 0);
  assign w595[26] = |(datain[207:204] ^ 15);
  assign w595[27] = |(datain[203:200] ^ 12);
  assign w595[28] = |(datain[199:196] ^ 7);
  assign w595[29] = |(datain[195:192] ^ 5);
  assign w595[30] = |(datain[191:188] ^ 0);
  assign w595[31] = |(datain[187:184] ^ 3);
  assign w595[32] = |(datain[183:180] ^ 14);
  assign w595[33] = |(datain[179:176] ^ 11);
  assign w595[34] = |(datain[175:172] ^ 5);
  assign w595[35] = |(datain[171:168] ^ 8);
  assign w595[36] = |(datain[167:164] ^ 9);
  assign w595[37] = |(datain[163:160] ^ 0);
  assign w595[38] = |(datain[159:156] ^ 15);
  assign w595[39] = |(datain[155:152] ^ 10);
  assign comp[595] = ~(|w595);
  wire [42-1:0] w596;
  assign w596[0] = |(datain[311:308] ^ 8);
  assign w596[1] = |(datain[307:304] ^ 11);
  assign w596[2] = |(datain[303:300] ^ 8);
  assign w596[3] = |(datain[299:296] ^ 11);
  assign w596[4] = |(datain[295:292] ^ 15);
  assign w596[5] = |(datain[291:288] ^ 2);
  assign w596[6] = |(datain[287:284] ^ 8);
  assign w596[7] = |(datain[283:280] ^ 11);
  assign w596[8] = |(datain[279:276] ^ 0);
  assign w596[9] = |(datain[275:272] ^ 4);
  assign w596[10] = |(datain[271:268] ^ 3);
  assign w596[11] = |(datain[267:264] ^ 2);
  assign w596[12] = |(datain[263:260] ^ 12);
  assign w596[13] = |(datain[259:256] ^ 4);
  assign w596[14] = |(datain[255:252] ^ 3);
  assign w596[15] = |(datain[251:248] ^ 12);
  assign w596[16] = |(datain[247:244] ^ 1);
  assign w596[17] = |(datain[243:240] ^ 7);
  assign w596[18] = |(datain[239:236] ^ 7);
  assign w596[19] = |(datain[235:232] ^ 4);
  assign w596[20] = |(datain[231:228] ^ 0);
  assign w596[21] = |(datain[227:224] ^ 11);
  assign w596[22] = |(datain[223:220] ^ 11);
  assign w596[23] = |(datain[219:216] ^ 8);
  assign w596[24] = |(datain[215:212] ^ 0);
  assign w596[25] = |(datain[211:208] ^ 0);
  assign w596[26] = |(datain[207:204] ^ 5);
  assign w596[27] = |(datain[203:200] ^ 7);
  assign w596[28] = |(datain[199:196] ^ 12);
  assign w596[29] = |(datain[195:192] ^ 13);
  assign w596[30] = |(datain[191:188] ^ 8);
  assign w596[31] = |(datain[187:184] ^ 11);
  assign w596[32] = |(datain[183:180] ^ 8);
  assign w596[33] = |(datain[179:176] ^ 3);
  assign w596[34] = |(datain[175:172] ^ 15);
  assign w596[35] = |(datain[171:168] ^ 1);
  assign w596[36] = |(datain[167:164] ^ 1);
  assign w596[37] = |(datain[163:160] ^ 15);
  assign w596[38] = |(datain[159:156] ^ 15);
  assign w596[39] = |(datain[155:152] ^ 6);
  assign w596[40] = |(datain[151:148] ^ 12);
  assign w596[41] = |(datain[147:144] ^ 1);
  assign comp[596] = ~(|w596);
  wire [76-1:0] w597;
  assign w597[0] = |(datain[311:308] ^ 15);
  assign w597[1] = |(datain[307:304] ^ 15);
  assign w597[2] = |(datain[303:300] ^ 4);
  assign w597[3] = |(datain[299:296] ^ 5);
  assign w597[4] = |(datain[295:292] ^ 4);
  assign w597[5] = |(datain[291:288] ^ 5);
  assign w597[6] = |(datain[287:284] ^ 12);
  assign w597[7] = |(datain[283:280] ^ 4);
  assign w597[8] = |(datain[279:276] ^ 3);
  assign w597[9] = |(datain[275:272] ^ 14);
  assign w597[10] = |(datain[271:268] ^ 8);
  assign w597[11] = |(datain[267:264] ^ 1);
  assign w597[12] = |(datain[263:260] ^ 0);
  assign w597[13] = |(datain[259:256] ^ 7);
  assign w597[14] = |(datain[255:252] ^ 2);
  assign w597[15] = |(datain[251:248] ^ 6);
  assign w597[16] = |(datain[247:244] ^ 8);
  assign w597[17] = |(datain[243:240] ^ 11);
  assign w597[18] = |(datain[239:236] ^ 7);
  assign w597[19] = |(datain[235:232] ^ 11);
  assign w597[20] = |(datain[231:228] ^ 7);
  assign w597[21] = |(datain[227:224] ^ 14);
  assign w597[22] = |(datain[223:220] ^ 10);
  assign w597[23] = |(datain[219:216] ^ 4);
  assign w597[24] = |(datain[215:212] ^ 10);
  assign w597[25] = |(datain[211:208] ^ 5);
  assign w597[26] = |(datain[207:204] ^ 7);
  assign w597[27] = |(datain[203:200] ^ 5);
  assign w597[28] = |(datain[199:196] ^ 15);
  assign w597[29] = |(datain[195:192] ^ 2);
  assign w597[30] = |(datain[191:188] ^ 1);
  assign w597[31] = |(datain[187:184] ^ 15);
  assign w597[32] = |(datain[183:180] ^ 5);
  assign w597[33] = |(datain[179:176] ^ 13);
  assign w597[34] = |(datain[175:172] ^ 5);
  assign w597[35] = |(datain[171:168] ^ 8);
  assign w597[36] = |(datain[167:164] ^ 2);
  assign w597[37] = |(datain[163:160] ^ 14);
  assign w597[38] = |(datain[159:156] ^ 15);
  assign w597[39] = |(datain[155:152] ^ 15);
  assign w597[40] = |(datain[151:148] ^ 3);
  assign w597[41] = |(datain[147:144] ^ 6);
  assign w597[42] = |(datain[143:140] ^ 8);
  assign w597[43] = |(datain[139:136] ^ 3);
  assign w597[44] = |(datain[135:132] ^ 0);
  assign w597[45] = |(datain[131:128] ^ 7);
  assign w597[46] = |(datain[127:124] ^ 5);
  assign w597[47] = |(datain[123:120] ^ 0);
  assign w597[48] = |(datain[119:116] ^ 5);
  assign w597[49] = |(datain[115:112] ^ 3);
  assign w597[50] = |(datain[111:108] ^ 11);
  assign w597[51] = |(datain[107:104] ^ 8);
  assign w597[52] = |(datain[103:100] ^ 2);
  assign w597[53] = |(datain[99:96] ^ 0);
  assign w597[54] = |(datain[95:92] ^ 1);
  assign w597[55] = |(datain[91:88] ^ 2);
  assign w597[56] = |(datain[87:84] ^ 12);
  assign w597[57] = |(datain[83:80] ^ 13);
  assign w597[58] = |(datain[79:76] ^ 2);
  assign w597[59] = |(datain[75:72] ^ 15);
  assign w597[60] = |(datain[71:68] ^ 2);
  assign w597[61] = |(datain[67:64] ^ 6);
  assign w597[62] = |(datain[63:60] ^ 8);
  assign w597[63] = |(datain[59:56] ^ 10);
  assign w597[64] = |(datain[55:52] ^ 1);
  assign w597[65] = |(datain[51:48] ^ 13);
  assign w597[66] = |(datain[47:44] ^ 11);
  assign w597[67] = |(datain[43:40] ^ 8);
  assign w597[68] = |(datain[39:36] ^ 1);
  assign w597[69] = |(datain[35:32] ^ 6);
  assign w597[70] = |(datain[31:28] ^ 1);
  assign w597[71] = |(datain[27:24] ^ 2);
  assign w597[72] = |(datain[23:20] ^ 12);
  assign w597[73] = |(datain[19:16] ^ 13);
  assign w597[74] = |(datain[15:12] ^ 2);
  assign w597[75] = |(datain[11:8] ^ 15);
  assign comp[597] = ~(|w597);
  wire [76-1:0] w598;
  assign w598[0] = |(datain[311:308] ^ 15);
  assign w598[1] = |(datain[307:304] ^ 15);
  assign w598[2] = |(datain[303:300] ^ 4);
  assign w598[3] = |(datain[299:296] ^ 5);
  assign w598[4] = |(datain[295:292] ^ 4);
  assign w598[5] = |(datain[291:288] ^ 5);
  assign w598[6] = |(datain[287:284] ^ 12);
  assign w598[7] = |(datain[283:280] ^ 4);
  assign w598[8] = |(datain[279:276] ^ 3);
  assign w598[9] = |(datain[275:272] ^ 14);
  assign w598[10] = |(datain[271:268] ^ 8);
  assign w598[11] = |(datain[267:264] ^ 15);
  assign w598[12] = |(datain[263:260] ^ 0);
  assign w598[13] = |(datain[259:256] ^ 7);
  assign w598[14] = |(datain[255:252] ^ 2);
  assign w598[15] = |(datain[251:248] ^ 6);
  assign w598[16] = |(datain[247:244] ^ 8);
  assign w598[17] = |(datain[243:240] ^ 11);
  assign w598[18] = |(datain[239:236] ^ 7);
  assign w598[19] = |(datain[235:232] ^ 11);
  assign w598[20] = |(datain[231:228] ^ 7);
  assign w598[21] = |(datain[227:224] ^ 14);
  assign w598[22] = |(datain[223:220] ^ 10);
  assign w598[23] = |(datain[219:216] ^ 4);
  assign w598[24] = |(datain[215:212] ^ 10);
  assign w598[25] = |(datain[211:208] ^ 5);
  assign w598[26] = |(datain[207:204] ^ 7);
  assign w598[27] = |(datain[203:200] ^ 5);
  assign w598[28] = |(datain[199:196] ^ 15);
  assign w598[29] = |(datain[195:192] ^ 2);
  assign w598[30] = |(datain[191:188] ^ 1);
  assign w598[31] = |(datain[187:184] ^ 15);
  assign w598[32] = |(datain[183:180] ^ 5);
  assign w598[33] = |(datain[179:176] ^ 13);
  assign w598[34] = |(datain[175:172] ^ 5);
  assign w598[35] = |(datain[171:168] ^ 8);
  assign w598[36] = |(datain[167:164] ^ 0);
  assign w598[37] = |(datain[163:160] ^ 6);
  assign w598[38] = |(datain[159:156] ^ 5);
  assign w598[39] = |(datain[155:152] ^ 0);
  assign w598[40] = |(datain[151:148] ^ 5);
  assign w598[41] = |(datain[147:144] ^ 3);
  assign w598[42] = |(datain[143:140] ^ 11);
  assign w598[43] = |(datain[139:136] ^ 8);
  assign w598[44] = |(datain[135:132] ^ 2);
  assign w598[45] = |(datain[131:128] ^ 0);
  assign w598[46] = |(datain[127:124] ^ 1);
  assign w598[47] = |(datain[123:120] ^ 2);
  assign w598[48] = |(datain[119:116] ^ 12);
  assign w598[49] = |(datain[115:112] ^ 13);
  assign w598[50] = |(datain[111:108] ^ 2);
  assign w598[51] = |(datain[107:104] ^ 15);
  assign w598[52] = |(datain[103:100] ^ 2);
  assign w598[53] = |(datain[99:96] ^ 6);
  assign w598[54] = |(datain[95:92] ^ 8);
  assign w598[55] = |(datain[91:88] ^ 10);
  assign w598[56] = |(datain[87:84] ^ 1);
  assign w598[57] = |(datain[83:80] ^ 13);
  assign w598[58] = |(datain[79:76] ^ 11);
  assign w598[59] = |(datain[75:72] ^ 8);
  assign w598[60] = |(datain[71:68] ^ 1);
  assign w598[61] = |(datain[67:64] ^ 6);
  assign w598[62] = |(datain[63:60] ^ 1);
  assign w598[63] = |(datain[59:56] ^ 2);
  assign w598[64] = |(datain[55:52] ^ 12);
  assign w598[65] = |(datain[51:48] ^ 13);
  assign w598[66] = |(datain[47:44] ^ 2);
  assign w598[67] = |(datain[43:40] ^ 15);
  assign w598[68] = |(datain[39:36] ^ 5);
  assign w598[69] = |(datain[35:32] ^ 11);
  assign w598[70] = |(datain[31:28] ^ 15);
  assign w598[71] = |(datain[27:24] ^ 15);
  assign w598[72] = |(datain[23:20] ^ 14);
  assign w598[73] = |(datain[19:16] ^ 5);
  assign w598[74] = |(datain[15:12] ^ 11);
  assign w598[75] = |(datain[11:8] ^ 14);
  assign comp[598] = ~(|w598);
  wire [40-1:0] w599;
  assign w599[0] = |(datain[311:308] ^ 15);
  assign w599[1] = |(datain[307:304] ^ 15);
  assign w599[2] = |(datain[303:300] ^ 11);
  assign w599[3] = |(datain[299:296] ^ 11);
  assign w599[4] = |(datain[295:292] ^ 1);
  assign w599[5] = |(datain[291:288] ^ 14);
  assign w599[6] = |(datain[287:284] ^ 0);
  assign w599[7] = |(datain[283:280] ^ 0);
  assign w599[8] = |(datain[279:276] ^ 11);
  assign w599[9] = |(datain[275:272] ^ 9);
  assign w599[10] = |(datain[271:268] ^ 12);
  assign w599[11] = |(datain[267:264] ^ 9);
  assign w599[12] = |(datain[263:260] ^ 1);
  assign w599[13] = |(datain[259:256] ^ 2);
  assign w599[14] = |(datain[255:252] ^ 0);
  assign w599[15] = |(datain[251:248] ^ 14);
  assign w599[16] = |(datain[247:244] ^ 1);
  assign w599[17] = |(datain[243:240] ^ 15);
  assign w599[18] = |(datain[239:236] ^ 13);
  assign w599[19] = |(datain[235:232] ^ 1);
  assign w599[20] = |(datain[231:228] ^ 14);
  assign w599[21] = |(datain[227:224] ^ 9);
  assign w599[22] = |(datain[223:220] ^ 8);
  assign w599[23] = |(datain[219:216] ^ 1);
  assign w599[24] = |(datain[215:212] ^ 3);
  assign w599[25] = |(datain[211:208] ^ 7);
  assign w599[26] = |(datain[207:204] ^ 1);
  assign w599[27] = |(datain[203:200] ^ 9);
  assign w599[28] = |(datain[199:196] ^ 3);
  assign w599[29] = |(datain[195:192] ^ 7);
  assign w599[30] = |(datain[191:188] ^ 8);
  assign w599[31] = |(datain[187:184] ^ 3);
  assign w599[32] = |(datain[183:180] ^ 12);
  assign w599[33] = |(datain[179:176] ^ 3);
  assign w599[34] = |(datain[175:172] ^ 0);
  assign w599[35] = |(datain[171:168] ^ 2);
  assign w599[36] = |(datain[167:164] ^ 14);
  assign w599[37] = |(datain[163:160] ^ 2);
  assign w599[38] = |(datain[159:156] ^ 15);
  assign w599[39] = |(datain[155:152] ^ 7);
  assign comp[599] = ~(|w599);
  wire [46-1:0] w600;
  assign w600[0] = |(datain[311:308] ^ 11);
  assign w600[1] = |(datain[307:304] ^ 8);
  assign w600[2] = |(datain[303:300] ^ 4);
  assign w600[3] = |(datain[299:296] ^ 4);
  assign w600[4] = |(datain[295:292] ^ 4);
  assign w600[5] = |(datain[291:288] ^ 1);
  assign w600[6] = |(datain[287:284] ^ 4);
  assign w600[7] = |(datain[283:280] ^ 12);
  assign w600[8] = |(datain[279:276] ^ 5);
  assign w600[9] = |(datain[275:272] ^ 6);
  assign w600[10] = |(datain[271:268] ^ 12);
  assign w600[11] = |(datain[267:264] ^ 13);
  assign w600[12] = |(datain[263:260] ^ 2);
  assign w600[13] = |(datain[259:256] ^ 1);
  assign w600[14] = |(datain[255:252] ^ 6);
  assign w600[15] = |(datain[251:248] ^ 6);
  assign w600[16] = |(datain[247:244] ^ 3);
  assign w600[17] = |(datain[243:240] ^ 13);
  assign w600[18] = |(datain[239:236] ^ 4);
  assign w600[19] = |(datain[235:232] ^ 11);
  assign w600[20] = |(datain[231:228] ^ 4);
  assign w600[21] = |(datain[227:224] ^ 3);
  assign w600[22] = |(datain[223:220] ^ 4);
  assign w600[23] = |(datain[219:216] ^ 15);
  assign w600[24] = |(datain[215:212] ^ 5);
  assign w600[25] = |(datain[211:208] ^ 2);
  assign w600[26] = |(datain[207:204] ^ 7);
  assign w600[27] = |(datain[203:200] ^ 4);
  assign w600[28] = |(datain[199:196] ^ 13);
  assign w600[29] = |(datain[195:192] ^ 5);
  assign w600[30] = |(datain[191:188] ^ 8);
  assign w600[31] = |(datain[187:184] ^ 12);
  assign w600[32] = |(datain[183:180] ^ 13);
  assign w600[33] = |(datain[179:176] ^ 8);
  assign w600[34] = |(datain[175:172] ^ 4);
  assign w600[35] = |(datain[171:168] ^ 8);
  assign w600[36] = |(datain[167:164] ^ 8);
  assign w600[37] = |(datain[163:160] ^ 14);
  assign w600[38] = |(datain[159:156] ^ 13);
  assign w600[39] = |(datain[155:152] ^ 8);
  assign w600[40] = |(datain[151:148] ^ 6);
  assign w600[41] = |(datain[147:144] ^ 6);
  assign w600[42] = |(datain[143:140] ^ 3);
  assign w600[43] = |(datain[139:136] ^ 3);
  assign w600[44] = |(datain[135:132] ^ 15);
  assign w600[45] = |(datain[131:128] ^ 15);
  assign comp[600] = ~(|w600);
  wire [74-1:0] w601;
  assign w601[0] = |(datain[311:308] ^ 1);
  assign w601[1] = |(datain[307:304] ^ 6);
  assign w601[2] = |(datain[303:300] ^ 8);
  assign w601[3] = |(datain[299:296] ^ 9);
  assign w601[4] = |(datain[295:292] ^ 1);
  assign w601[5] = |(datain[291:288] ^ 6);
  assign w601[6] = |(datain[287:284] ^ 0);
  assign w601[7] = |(datain[283:280] ^ 1);
  assign w601[8] = |(datain[279:276] ^ 0);
  assign w601[9] = |(datain[275:272] ^ 0);
  assign w601[10] = |(datain[271:268] ^ 8);
  assign w601[11] = |(datain[267:264] ^ 1);
  assign w601[12] = |(datain[263:260] ^ 12);
  assign w601[13] = |(datain[259:256] ^ 2);
  assign w601[14] = |(datain[255:252] ^ 10);
  assign w601[15] = |(datain[251:248] ^ 2);
  assign w601[16] = |(datain[247:244] ^ 0);
  assign w601[17] = |(datain[243:240] ^ 4);
  assign w601[18] = |(datain[239:236] ^ 8);
  assign w601[19] = |(datain[235:232] ^ 3);
  assign w601[20] = |(datain[231:228] ^ 14);
  assign w601[21] = |(datain[227:224] ^ 2);
  assign w601[22] = |(datain[223:220] ^ 15);
  assign w601[23] = |(datain[219:216] ^ 14);
  assign w601[24] = |(datain[215:212] ^ 4);
  assign w601[25] = |(datain[211:208] ^ 0);
  assign w601[26] = |(datain[207:204] ^ 6);
  assign w601[27] = |(datain[203:200] ^ 7);
  assign w601[28] = |(datain[199:196] ^ 8);
  assign w601[29] = |(datain[195:192] ^ 9);
  assign w601[30] = |(datain[191:188] ^ 4);
  assign w601[31] = |(datain[187:184] ^ 6);
  assign w601[32] = |(datain[183:180] ^ 0);
  assign w601[33] = |(datain[179:176] ^ 14);
  assign w601[34] = |(datain[175:172] ^ 6);
  assign w601[35] = |(datain[171:168] ^ 7);
  assign w601[36] = |(datain[167:164] ^ 8);
  assign w601[37] = |(datain[163:160] ^ 9);
  assign w601[38] = |(datain[159:156] ^ 5);
  assign w601[39] = |(datain[155:152] ^ 6);
  assign w601[40] = |(datain[151:148] ^ 1);
  assign w601[41] = |(datain[147:144] ^ 0);
  assign w601[42] = |(datain[143:140] ^ 11);
  assign w601[43] = |(datain[139:136] ^ 4);
  assign w601[44] = |(datain[135:132] ^ 4);
  assign w601[45] = |(datain[131:128] ^ 0);
  assign w601[46] = |(datain[127:124] ^ 11);
  assign w601[47] = |(datain[123:120] ^ 9);
  assign w601[48] = |(datain[119:116] ^ 8);
  assign w601[49] = |(datain[115:112] ^ 13);
  assign w601[50] = |(datain[111:108] ^ 0);
  assign w601[51] = |(datain[107:104] ^ 2);
  assign w601[52] = |(datain[103:100] ^ 3);
  assign w601[53] = |(datain[99:96] ^ 3);
  assign w601[54] = |(datain[95:92] ^ 13);
  assign w601[55] = |(datain[91:88] ^ 2);
  assign w601[56] = |(datain[87:84] ^ 14);
  assign w601[57] = |(datain[83:80] ^ 8);
  assign w601[58] = |(datain[79:76] ^ 5);
  assign w601[59] = |(datain[75:72] ^ 15);
  assign w601[60] = |(datain[71:68] ^ 15);
  assign w601[61] = |(datain[67:64] ^ 15);
  assign w601[62] = |(datain[63:60] ^ 14);
  assign w601[63] = |(datain[59:56] ^ 8);
  assign w601[64] = |(datain[55:52] ^ 3);
  assign w601[65] = |(datain[51:48] ^ 6);
  assign w601[66] = |(datain[47:44] ^ 0);
  assign w601[67] = |(datain[43:40] ^ 0);
  assign w601[68] = |(datain[39:36] ^ 11);
  assign w601[69] = |(datain[35:32] ^ 9);
  assign w601[70] = |(datain[31:28] ^ 0);
  assign w601[71] = |(datain[27:24] ^ 0);
  assign w601[72] = |(datain[23:20] ^ 0);
  assign w601[73] = |(datain[19:16] ^ 2);
  assign comp[601] = ~(|w601);
  wire [30-1:0] w602;
  assign w602[0] = |(datain[311:308] ^ 14);
  assign w602[1] = |(datain[307:304] ^ 2);
  assign w602[2] = |(datain[303:300] ^ 0);
  assign w602[3] = |(datain[299:296] ^ 1);
  assign w602[4] = |(datain[295:292] ^ 11);
  assign w602[5] = |(datain[291:288] ^ 10);
  assign w602[6] = |(datain[287:284] ^ 7);
  assign w602[7] = |(datain[283:280] ^ 0);
  assign w602[8] = |(datain[279:276] ^ 0);
  assign w602[9] = |(datain[275:272] ^ 1);
  assign w602[10] = |(datain[271:268] ^ 2);
  assign w602[11] = |(datain[267:264] ^ 14);
  assign w602[12] = |(datain[263:260] ^ 8);
  assign w602[13] = |(datain[259:256] ^ 1);
  assign w602[14] = |(datain[255:252] ^ 3);
  assign w602[15] = |(datain[251:248] ^ 4);
  assign w602[16] = |(datain[247:244] ^ 2);
  assign w602[17] = |(datain[243:240] ^ 8);
  assign w602[18] = |(datain[239:236] ^ 3);
  assign w602[19] = |(datain[235:232] ^ 1);
  assign w602[20] = |(datain[231:228] ^ 4);
  assign w602[21] = |(datain[227:224] ^ 6);
  assign w602[22] = |(datain[223:220] ^ 4);
  assign w602[23] = |(datain[219:216] ^ 6);
  assign w602[24] = |(datain[215:212] ^ 4);
  assign w602[25] = |(datain[211:208] ^ 10);
  assign w602[26] = |(datain[207:204] ^ 7);
  assign w602[27] = |(datain[203:200] ^ 5);
  assign w602[28] = |(datain[199:196] ^ 15);
  assign w602[29] = |(datain[195:192] ^ 6);
  assign comp[602] = ~(|w602);
  wire [74-1:0] w603;
  assign w603[0] = |(datain[311:308] ^ 5);
  assign w603[1] = |(datain[307:304] ^ 3);
  assign w603[2] = |(datain[303:300] ^ 5);
  assign w603[3] = |(datain[299:296] ^ 6);
  assign w603[4] = |(datain[295:292] ^ 5);
  assign w603[5] = |(datain[291:288] ^ 7);
  assign w603[6] = |(datain[287:284] ^ 15);
  assign w603[7] = |(datain[283:280] ^ 10);
  assign w603[8] = |(datain[279:276] ^ 8);
  assign w603[9] = |(datain[275:272] ^ 12);
  assign w603[10] = |(datain[271:268] ^ 12);
  assign w603[11] = |(datain[267:264] ^ 8);
  assign w603[12] = |(datain[263:260] ^ 8);
  assign w603[13] = |(datain[259:256] ^ 14);
  assign w603[14] = |(datain[255:252] ^ 13);
  assign w603[15] = |(datain[251:248] ^ 8);
  assign w603[16] = |(datain[247:244] ^ 8);
  assign w603[17] = |(datain[243:240] ^ 14);
  assign w603[18] = |(datain[239:236] ^ 12);
  assign w603[19] = |(datain[235:232] ^ 0);
  assign w603[20] = |(datain[231:228] ^ 11);
  assign w603[21] = |(datain[227:224] ^ 14);
  assign w603[22] = |(datain[223:220] ^ 7);
  assign w603[23] = |(datain[219:216] ^ 8);
  assign w603[24] = |(datain[215:212] ^ 0);
  assign w603[25] = |(datain[211:208] ^ 0);
  assign w603[26] = |(datain[207:204] ^ 0);
  assign w603[27] = |(datain[203:200] ^ 3);
  assign w603[28] = |(datain[199:196] ^ 15);
  assign w603[29] = |(datain[195:192] ^ 5);
  assign w603[30] = |(datain[191:188] ^ 8);
  assign w603[31] = |(datain[187:184] ^ 11);
  assign w603[32] = |(datain[183:180] ^ 15);
  assign w603[33] = |(datain[179:176] ^ 14);
  assign w603[34] = |(datain[175:172] ^ 11);
  assign w603[35] = |(datain[171:168] ^ 9);
  assign w603[36] = |(datain[167:164] ^ 8);
  assign w603[37] = |(datain[163:160] ^ 11);
  assign w603[38] = |(datain[159:156] ^ 0);
  assign w603[39] = |(datain[155:152] ^ 1);
  assign w603[40] = |(datain[151:148] ^ 8);
  assign w603[41] = |(datain[147:144] ^ 11);
  assign w603[42] = |(datain[143:140] ^ 13);
  assign w603[43] = |(datain[139:136] ^ 13);
  assign w603[44] = |(datain[135:132] ^ 15);
  assign w603[45] = |(datain[131:128] ^ 12);
  assign w603[46] = |(datain[127:124] ^ 10);
  assign w603[47] = |(datain[123:120] ^ 13);
  assign w603[48] = |(datain[119:116] ^ 3);
  assign w603[49] = |(datain[115:112] ^ 3);
  assign w603[50] = |(datain[111:108] ^ 8);
  assign w603[51] = |(datain[107:104] ^ 7);
  assign w603[52] = |(datain[103:100] ^ 6);
  assign w603[53] = |(datain[99:96] ^ 0);
  assign w603[54] = |(datain[95:92] ^ 0);
  assign w603[55] = |(datain[91:88] ^ 0);
  assign w603[56] = |(datain[87:84] ^ 10);
  assign w603[57] = |(datain[83:80] ^ 11);
  assign w603[58] = |(datain[79:76] ^ 14);
  assign w603[59] = |(datain[75:72] ^ 2);
  assign w603[60] = |(datain[71:68] ^ 15);
  assign w603[61] = |(datain[67:64] ^ 8);
  assign w603[62] = |(datain[63:60] ^ 5);
  assign w603[63] = |(datain[59:56] ^ 15);
  assign w603[64] = |(datain[55:52] ^ 5);
  assign w603[65] = |(datain[51:48] ^ 14);
  assign w603[66] = |(datain[47:44] ^ 5);
  assign w603[67] = |(datain[43:40] ^ 11);
  assign w603[68] = |(datain[39:36] ^ 0);
  assign w603[69] = |(datain[35:32] ^ 7);
  assign w603[70] = |(datain[31:28] ^ 1);
  assign w603[71] = |(datain[27:24] ^ 15);
  assign w603[72] = |(datain[23:20] ^ 12);
  assign w603[73] = |(datain[19:16] ^ 3);
  assign comp[603] = ~(|w603);
  wire [74-1:0] w604;
  assign w604[0] = |(datain[311:308] ^ 13);
  assign w604[1] = |(datain[307:304] ^ 8);
  assign w604[2] = |(datain[303:300] ^ 10);
  assign w604[3] = |(datain[299:296] ^ 1);
  assign w604[4] = |(datain[295:292] ^ 8);
  assign w604[5] = |(datain[291:288] ^ 4);
  assign w604[6] = |(datain[287:284] ^ 0);
  assign w604[7] = |(datain[283:280] ^ 0);
  assign w604[8] = |(datain[279:276] ^ 2);
  assign w604[9] = |(datain[275:272] ^ 14);
  assign w604[10] = |(datain[271:268] ^ 10);
  assign w604[11] = |(datain[267:264] ^ 3);
  assign w604[12] = |(datain[263:260] ^ 12);
  assign w604[13] = |(datain[259:256] ^ 13);
  assign w604[14] = |(datain[255:252] ^ 0);
  assign w604[15] = |(datain[251:248] ^ 1);
  assign w604[16] = |(datain[247:244] ^ 10);
  assign w604[17] = |(datain[243:240] ^ 1);
  assign w604[18] = |(datain[239:236] ^ 8);
  assign w604[19] = |(datain[235:232] ^ 6);
  assign w604[20] = |(datain[231:228] ^ 0);
  assign w604[21] = |(datain[227:224] ^ 0);
  assign w604[22] = |(datain[223:220] ^ 2);
  assign w604[23] = |(datain[219:216] ^ 14);
  assign w604[24] = |(datain[215:212] ^ 10);
  assign w604[25] = |(datain[211:208] ^ 3);
  assign w604[26] = |(datain[207:204] ^ 12);
  assign w604[27] = |(datain[203:200] ^ 15);
  assign w604[28] = |(datain[199:196] ^ 0);
  assign w604[29] = |(datain[195:192] ^ 1);
  assign w604[30] = |(datain[191:188] ^ 11);
  assign w604[31] = |(datain[187:184] ^ 8);
  assign w604[32] = |(datain[183:180] ^ 0);
  assign w604[33] = |(datain[179:176] ^ 5);
  assign w604[34] = |(datain[175:172] ^ 15);
  assign w604[35] = |(datain[171:168] ^ 15);
  assign w604[36] = |(datain[167:164] ^ 9);
  assign w604[37] = |(datain[163:160] ^ 12);
  assign w604[38] = |(datain[159:156] ^ 2);
  assign w604[39] = |(datain[155:152] ^ 14);
  assign w604[40] = |(datain[151:148] ^ 15);
  assign w604[41] = |(datain[147:144] ^ 15);
  assign w604[42] = |(datain[143:140] ^ 1);
  assign w604[43] = |(datain[139:136] ^ 14);
  assign w604[44] = |(datain[135:132] ^ 12);
  assign w604[45] = |(datain[131:128] ^ 13);
  assign w604[46] = |(datain[127:124] ^ 0);
  assign w604[47] = |(datain[123:120] ^ 1);
  assign w604[48] = |(datain[119:116] ^ 3);
  assign w604[49] = |(datain[115:112] ^ 13);
  assign w604[50] = |(datain[111:108] ^ 15);
  assign w604[51] = |(datain[107:104] ^ 15);
  assign w604[52] = |(datain[103:100] ^ 0);
  assign w604[53] = |(datain[99:96] ^ 5);
  assign w604[54] = |(datain[95:92] ^ 7);
  assign w604[55] = |(datain[91:88] ^ 4);
  assign w604[56] = |(datain[87:84] ^ 1);
  assign w604[57] = |(datain[83:80] ^ 14);
  assign w604[58] = |(datain[79:76] ^ 15);
  assign w604[59] = |(datain[75:72] ^ 12);
  assign w604[60] = |(datain[71:68] ^ 3);
  assign w604[61] = |(datain[67:64] ^ 3);
  assign w604[62] = |(datain[63:60] ^ 15);
  assign w604[63] = |(datain[59:56] ^ 6);
  assign w604[64] = |(datain[55:52] ^ 8);
  assign w604[65] = |(datain[51:48] ^ 14);
  assign w604[66] = |(datain[47:44] ^ 12);
  assign w604[67] = |(datain[43:40] ^ 6);
  assign w604[68] = |(datain[39:36] ^ 0);
  assign w604[69] = |(datain[35:32] ^ 14);
  assign w604[70] = |(datain[31:28] ^ 1);
  assign w604[71] = |(datain[27:24] ^ 15);
  assign w604[72] = |(datain[23:20] ^ 11);
  assign w604[73] = |(datain[19:16] ^ 15);
  assign comp[604] = ~(|w604);
  wire [72-1:0] w605;
  assign w605[0] = |(datain[311:308] ^ 0);
  assign w605[1] = |(datain[307:304] ^ 2);
  assign w605[2] = |(datain[303:300] ^ 0);
  assign w605[3] = |(datain[299:296] ^ 0);
  assign w605[4] = |(datain[295:292] ^ 11);
  assign w605[5] = |(datain[291:288] ^ 4);
  assign w605[6] = |(datain[287:284] ^ 4);
  assign w605[7] = |(datain[283:280] ^ 0);
  assign w605[8] = |(datain[279:276] ^ 9);
  assign w605[9] = |(datain[275:272] ^ 12);
  assign w605[10] = |(datain[271:268] ^ 2);
  assign w605[11] = |(datain[267:264] ^ 14);
  assign w605[12] = |(datain[263:260] ^ 15);
  assign w605[13] = |(datain[259:256] ^ 15);
  assign w605[14] = |(datain[255:252] ^ 1);
  assign w605[15] = |(datain[251:248] ^ 14);
  assign w605[16] = |(datain[247:244] ^ 12);
  assign w605[17] = |(datain[243:240] ^ 13);
  assign w605[18] = |(datain[239:236] ^ 0);
  assign w605[19] = |(datain[235:232] ^ 0);
  assign w605[20] = |(datain[231:228] ^ 3);
  assign w605[21] = |(datain[227:224] ^ 3);
  assign w605[22] = |(datain[223:220] ^ 12);
  assign w605[23] = |(datain[219:216] ^ 9);
  assign w605[24] = |(datain[215:212] ^ 8);
  assign w605[25] = |(datain[211:208] ^ 11);
  assign w605[26] = |(datain[207:204] ^ 1);
  assign w605[27] = |(datain[203:200] ^ 6);
  assign w605[28] = |(datain[199:196] ^ 1);
  assign w605[29] = |(datain[195:192] ^ 6);
  assign w605[30] = |(datain[191:188] ^ 0);
  assign w605[31] = |(datain[187:184] ^ 0);
  assign w605[32] = |(datain[183:180] ^ 8);
  assign w605[33] = |(datain[179:176] ^ 1);
  assign w605[34] = |(datain[175:172] ^ 12);
  assign w605[35] = |(datain[171:168] ^ 2);
  assign w605[36] = |(datain[167:164] ^ 8);
  assign w605[37] = |(datain[163:160] ^ 13);
  assign w605[38] = |(datain[159:156] ^ 1);
  assign w605[39] = |(datain[155:152] ^ 14);
  assign w605[40] = |(datain[151:148] ^ 11);
  assign w605[41] = |(datain[147:144] ^ 8);
  assign w605[42] = |(datain[143:140] ^ 0);
  assign w605[43] = |(datain[139:136] ^ 0);
  assign w605[44] = |(datain[135:132] ^ 4);
  assign w605[45] = |(datain[131:128] ^ 2);
  assign w605[46] = |(datain[127:124] ^ 9);
  assign w605[47] = |(datain[123:120] ^ 12);
  assign w605[48] = |(datain[119:116] ^ 2);
  assign w605[49] = |(datain[115:112] ^ 14);
  assign w605[50] = |(datain[111:108] ^ 15);
  assign w605[51] = |(datain[107:104] ^ 15);
  assign w605[52] = |(datain[103:100] ^ 1);
  assign w605[53] = |(datain[99:96] ^ 14);
  assign w605[54] = |(datain[95:92] ^ 12);
  assign w605[55] = |(datain[91:88] ^ 13);
  assign w605[56] = |(datain[87:84] ^ 0);
  assign w605[57] = |(datain[83:80] ^ 0);
  assign w605[58] = |(datain[79:76] ^ 11);
  assign w605[59] = |(datain[75:72] ^ 4);
  assign w605[60] = |(datain[71:68] ^ 4);
  assign w605[61] = |(datain[67:64] ^ 0);
  assign w605[62] = |(datain[63:60] ^ 9);
  assign w605[63] = |(datain[59:56] ^ 12);
  assign w605[64] = |(datain[55:52] ^ 2);
  assign w605[65] = |(datain[51:48] ^ 14);
  assign w605[66] = |(datain[47:44] ^ 15);
  assign w605[67] = |(datain[43:40] ^ 15);
  assign w605[68] = |(datain[39:36] ^ 1);
  assign w605[69] = |(datain[35:32] ^ 14);
  assign w605[70] = |(datain[31:28] ^ 12);
  assign w605[71] = |(datain[27:24] ^ 13);
  assign comp[605] = ~(|w605);
  wire [76-1:0] w606;
  assign w606[0] = |(datain[311:308] ^ 0);
  assign w606[1] = |(datain[307:304] ^ 6);
  assign w606[2] = |(datain[303:300] ^ 5);
  assign w606[3] = |(datain[299:296] ^ 3);
  assign w606[4] = |(datain[295:292] ^ 5);
  assign w606[5] = |(datain[291:288] ^ 6);
  assign w606[6] = |(datain[287:284] ^ 5);
  assign w606[7] = |(datain[283:280] ^ 7);
  assign w606[8] = |(datain[279:276] ^ 15);
  assign w606[9] = |(datain[275:272] ^ 10);
  assign w606[10] = |(datain[271:268] ^ 8);
  assign w606[11] = |(datain[267:264] ^ 12);
  assign w606[12] = |(datain[263:260] ^ 12);
  assign w606[13] = |(datain[259:256] ^ 8);
  assign w606[14] = |(datain[255:252] ^ 8);
  assign w606[15] = |(datain[251:248] ^ 14);
  assign w606[16] = |(datain[247:244] ^ 13);
  assign w606[17] = |(datain[243:240] ^ 8);
  assign w606[18] = |(datain[239:236] ^ 8);
  assign w606[19] = |(datain[235:232] ^ 14);
  assign w606[20] = |(datain[231:228] ^ 12);
  assign w606[21] = |(datain[227:224] ^ 0);
  assign w606[22] = |(datain[223:220] ^ 11);
  assign w606[23] = |(datain[219:216] ^ 14);
  assign w606[24] = |(datain[215:212] ^ 5);
  assign w606[25] = |(datain[211:208] ^ 14);
  assign w606[26] = |(datain[207:204] ^ 0);
  assign w606[27] = |(datain[203:200] ^ 0);
  assign w606[28] = |(datain[199:196] ^ 0);
  assign w606[29] = |(datain[195:192] ^ 3);
  assign w606[30] = |(datain[191:188] ^ 15);
  assign w606[31] = |(datain[187:184] ^ 5);
  assign w606[32] = |(datain[183:180] ^ 8);
  assign w606[33] = |(datain[179:176] ^ 11);
  assign w606[34] = |(datain[175:172] ^ 15);
  assign w606[35] = |(datain[171:168] ^ 14);
  assign w606[36] = |(datain[167:164] ^ 11);
  assign w606[37] = |(datain[163:160] ^ 9);
  assign w606[38] = |(datain[159:156] ^ 11);
  assign w606[39] = |(datain[155:152] ^ 1);
  assign w606[40] = |(datain[151:148] ^ 0);
  assign w606[41] = |(datain[147:144] ^ 2);
  assign w606[42] = |(datain[143:140] ^ 8);
  assign w606[43] = |(datain[139:136] ^ 11);
  assign w606[44] = |(datain[135:132] ^ 13);
  assign w606[45] = |(datain[131:128] ^ 13);
  assign w606[46] = |(datain[127:124] ^ 15);
  assign w606[47] = |(datain[123:120] ^ 12);
  assign w606[48] = |(datain[119:116] ^ 10);
  assign w606[49] = |(datain[115:112] ^ 13);
  assign w606[50] = |(datain[111:108] ^ 3);
  assign w606[51] = |(datain[107:104] ^ 3);
  assign w606[52] = |(datain[103:100] ^ 8);
  assign w606[53] = |(datain[99:96] ^ 7);
  assign w606[54] = |(datain[95:92] ^ 3);
  assign w606[55] = |(datain[91:88] ^ 15);
  assign w606[56] = |(datain[87:84] ^ 0);
  assign w606[57] = |(datain[83:80] ^ 0);
  assign w606[58] = |(datain[79:76] ^ 10);
  assign w606[59] = |(datain[75:72] ^ 11);
  assign w606[60] = |(datain[71:68] ^ 14);
  assign w606[61] = |(datain[67:64] ^ 2);
  assign w606[62] = |(datain[63:60] ^ 15);
  assign w606[63] = |(datain[59:56] ^ 8);
  assign w606[64] = |(datain[55:52] ^ 5);
  assign w606[65] = |(datain[51:48] ^ 15);
  assign w606[66] = |(datain[47:44] ^ 5);
  assign w606[67] = |(datain[43:40] ^ 14);
  assign w606[68] = |(datain[39:36] ^ 5);
  assign w606[69] = |(datain[35:32] ^ 11);
  assign w606[70] = |(datain[31:28] ^ 0);
  assign w606[71] = |(datain[27:24] ^ 7);
  assign w606[72] = |(datain[23:20] ^ 1);
  assign w606[73] = |(datain[19:16] ^ 15);
  assign w606[74] = |(datain[15:12] ^ 12);
  assign w606[75] = |(datain[11:8] ^ 3);
  assign comp[606] = ~(|w606);
  wire [46-1:0] w607;
  assign w607[0] = |(datain[311:308] ^ 8);
  assign w607[1] = |(datain[307:304] ^ 14);
  assign w607[2] = |(datain[303:300] ^ 12);
  assign w607[3] = |(datain[299:296] ^ 0);
  assign w607[4] = |(datain[295:292] ^ 11);
  assign w607[5] = |(datain[291:288] ^ 14);
  assign w607[6] = |(datain[287:284] ^ 7);
  assign w607[7] = |(datain[283:280] ^ 9);
  assign w607[8] = |(datain[279:276] ^ 0);
  assign w607[9] = |(datain[275:272] ^ 0);
  assign w607[10] = |(datain[271:268] ^ 0);
  assign w607[11] = |(datain[267:264] ^ 3);
  assign w607[12] = |(datain[263:260] ^ 15);
  assign w607[13] = |(datain[259:256] ^ 5);
  assign w607[14] = |(datain[255:252] ^ 8);
  assign w607[15] = |(datain[251:248] ^ 11);
  assign w607[16] = |(datain[247:244] ^ 15);
  assign w607[17] = |(datain[243:240] ^ 14);
  assign w607[18] = |(datain[239:236] ^ 11);
  assign w607[19] = |(datain[235:232] ^ 9);
  assign w607[20] = |(datain[231:228] ^ 6);
  assign w607[21] = |(datain[227:224] ^ 15);
  assign w607[22] = |(datain[223:220] ^ 0);
  assign w607[23] = |(datain[219:216] ^ 1);
  assign w607[24] = |(datain[215:212] ^ 8);
  assign w607[25] = |(datain[211:208] ^ 11);
  assign w607[26] = |(datain[207:204] ^ 13);
  assign w607[27] = |(datain[203:200] ^ 13);
  assign w607[28] = |(datain[199:196] ^ 15);
  assign w607[29] = |(datain[195:192] ^ 12);
  assign w607[30] = |(datain[191:188] ^ 10);
  assign w607[31] = |(datain[187:184] ^ 13);
  assign w607[32] = |(datain[183:180] ^ 3);
  assign w607[33] = |(datain[179:176] ^ 3);
  assign w607[34] = |(datain[175:172] ^ 8);
  assign w607[35] = |(datain[171:168] ^ 7);
  assign w607[36] = |(datain[167:164] ^ 6);
  assign w607[37] = |(datain[163:160] ^ 7);
  assign w607[38] = |(datain[159:156] ^ 0);
  assign w607[39] = |(datain[155:152] ^ 0);
  assign w607[40] = |(datain[151:148] ^ 10);
  assign w607[41] = |(datain[147:144] ^ 11);
  assign w607[42] = |(datain[143:140] ^ 14);
  assign w607[43] = |(datain[139:136] ^ 2);
  assign w607[44] = |(datain[135:132] ^ 15);
  assign w607[45] = |(datain[131:128] ^ 8);
  assign comp[607] = ~(|w607);
  wire [46-1:0] w608;
  assign w608[0] = |(datain[311:308] ^ 0);
  assign w608[1] = |(datain[307:304] ^ 11);
  assign w608[2] = |(datain[303:300] ^ 0);
  assign w608[3] = |(datain[299:296] ^ 0);
  assign w608[4] = |(datain[295:292] ^ 0);
  assign w608[5] = |(datain[291:288] ^ 3);
  assign w608[6] = |(datain[287:284] ^ 15);
  assign w608[7] = |(datain[283:280] ^ 5);
  assign w608[8] = |(datain[279:276] ^ 8);
  assign w608[9] = |(datain[275:272] ^ 11);
  assign w608[10] = |(datain[271:268] ^ 15);
  assign w608[11] = |(datain[267:264] ^ 14);
  assign w608[12] = |(datain[263:260] ^ 11);
  assign w608[13] = |(datain[259:256] ^ 9);
  assign w608[14] = |(datain[255:252] ^ 8);
  assign w608[15] = |(datain[251:248] ^ 4);
  assign w608[16] = |(datain[247:244] ^ 0);
  assign w608[17] = |(datain[243:240] ^ 1);
  assign w608[18] = |(datain[239:236] ^ 8);
  assign w608[19] = |(datain[235:232] ^ 11);
  assign w608[20] = |(datain[231:228] ^ 13);
  assign w608[21] = |(datain[227:224] ^ 13);
  assign w608[22] = |(datain[223:220] ^ 15);
  assign w608[23] = |(datain[219:216] ^ 12);
  assign w608[24] = |(datain[215:212] ^ 10);
  assign w608[25] = |(datain[211:208] ^ 13);
  assign w608[26] = |(datain[207:204] ^ 2);
  assign w608[27] = |(datain[203:200] ^ 14);
  assign w608[28] = |(datain[199:196] ^ 3);
  assign w608[29] = |(datain[195:192] ^ 3);
  assign w608[30] = |(datain[191:188] ^ 8);
  assign w608[31] = |(datain[187:184] ^ 7);
  assign w608[32] = |(datain[183:180] ^ 12);
  assign w608[33] = |(datain[179:176] ^ 11);
  assign w608[34] = |(datain[175:172] ^ 0);
  assign w608[35] = |(datain[171:168] ^ 3);
  assign w608[36] = |(datain[167:164] ^ 10);
  assign w608[37] = |(datain[163:160] ^ 11);
  assign w608[38] = |(datain[159:156] ^ 14);
  assign w608[39] = |(datain[155:152] ^ 2);
  assign w608[40] = |(datain[151:148] ^ 15);
  assign w608[41] = |(datain[147:144] ^ 7);
  assign w608[42] = |(datain[143:140] ^ 5);
  assign w608[43] = |(datain[139:136] ^ 11);
  assign w608[44] = |(datain[135:132] ^ 0);
  assign w608[45] = |(datain[131:128] ^ 7);
  assign comp[608] = ~(|w608);
  wire [42-1:0] w609;
  assign w609[0] = |(datain[311:308] ^ 2);
  assign w609[1] = |(datain[307:304] ^ 0);
  assign w609[2] = |(datain[303:300] ^ 0);
  assign w609[3] = |(datain[299:296] ^ 4);
  assign w609[4] = |(datain[295:292] ^ 11);
  assign w609[5] = |(datain[291:288] ^ 4);
  assign w609[6] = |(datain[287:284] ^ 4);
  assign w609[7] = |(datain[283:280] ^ 0);
  assign w609[8] = |(datain[279:276] ^ 12);
  assign w609[9] = |(datain[275:272] ^ 13);
  assign w609[10] = |(datain[271:268] ^ 2);
  assign w609[11] = |(datain[267:264] ^ 1);
  assign w609[12] = |(datain[263:260] ^ 11);
  assign w609[13] = |(datain[259:256] ^ 4);
  assign w609[14] = |(datain[255:252] ^ 3);
  assign w609[15] = |(datain[251:248] ^ 14);
  assign w609[16] = |(datain[247:244] ^ 12);
  assign w609[17] = |(datain[243:240] ^ 13);
  assign w609[18] = |(datain[239:236] ^ 2);
  assign w609[19] = |(datain[235:232] ^ 1);
  assign w609[20] = |(datain[231:228] ^ 5);
  assign w609[21] = |(datain[227:224] ^ 8);
  assign w609[22] = |(datain[223:220] ^ 8);
  assign w609[23] = |(datain[219:216] ^ 14);
  assign w609[24] = |(datain[215:212] ^ 13);
  assign w609[25] = |(datain[211:208] ^ 8);
  assign w609[26] = |(datain[207:204] ^ 5);
  assign w609[27] = |(datain[203:200] ^ 10);
  assign w609[28] = |(datain[199:196] ^ 11);
  assign w609[29] = |(datain[195:192] ^ 8);
  assign w609[30] = |(datain[191:188] ^ 0);
  assign w609[31] = |(datain[187:184] ^ 1);
  assign w609[32] = |(datain[183:180] ^ 4);
  assign w609[33] = |(datain[179:176] ^ 3);
  assign w609[34] = |(datain[175:172] ^ 11);
  assign w609[35] = |(datain[171:168] ^ 9);
  assign w609[36] = |(datain[167:164] ^ 0);
  assign w609[37] = |(datain[163:160] ^ 1);
  assign w609[38] = |(datain[159:156] ^ 0);
  assign w609[39] = |(datain[155:152] ^ 0);
  assign w609[40] = |(datain[151:148] ^ 12);
  assign w609[41] = |(datain[147:144] ^ 13);
  assign comp[609] = ~(|w609);
  wire [44-1:0] w610;
  assign w610[0] = |(datain[311:308] ^ 4);
  assign w610[1] = |(datain[307:304] ^ 2);
  assign w610[2] = |(datain[303:300] ^ 8);
  assign w610[3] = |(datain[299:296] ^ 11);
  assign w610[4] = |(datain[295:292] ^ 12);
  assign w610[5] = |(datain[291:288] ^ 10);
  assign w610[6] = |(datain[287:284] ^ 12);
  assign w610[7] = |(datain[283:280] ^ 13);
  assign w610[8] = |(datain[279:276] ^ 3);
  assign w610[9] = |(datain[275:272] ^ 5);
  assign w610[10] = |(datain[271:268] ^ 11);
  assign w610[11] = |(datain[267:264] ^ 4);
  assign w610[12] = |(datain[263:260] ^ 4);
  assign w610[13] = |(datain[259:256] ^ 0);
  assign w610[14] = |(datain[255:252] ^ 11);
  assign w610[15] = |(datain[251:248] ^ 2);
  assign w610[16] = |(datain[247:244] ^ 2);
  assign w610[17] = |(datain[243:240] ^ 13);
  assign w610[18] = |(datain[239:236] ^ 11);
  assign w610[19] = |(datain[235:232] ^ 1);
  assign w610[20] = |(datain[231:228] ^ 0);
  assign w610[21] = |(datain[227:224] ^ 3);
  assign w610[22] = |(datain[223:220] ^ 8);
  assign w610[23] = |(datain[219:216] ^ 9);
  assign w610[24] = |(datain[215:212] ^ 2);
  assign w610[25] = |(datain[211:208] ^ 12);
  assign w610[26] = |(datain[207:204] ^ 12);
  assign w610[27] = |(datain[203:200] ^ 13);
  assign w610[28] = |(datain[199:196] ^ 14);
  assign w610[29] = |(datain[195:192] ^ 5);
  assign w610[30] = |(datain[191:188] ^ 11);
  assign w610[31] = |(datain[187:184] ^ 4);
  assign w610[32] = |(datain[183:180] ^ 3);
  assign w610[33] = |(datain[179:176] ^ 14);
  assign w610[34] = |(datain[175:172] ^ 12);
  assign w610[35] = |(datain[171:168] ^ 13);
  assign w610[36] = |(datain[167:164] ^ 14);
  assign w610[37] = |(datain[163:160] ^ 5);
  assign w610[38] = |(datain[159:156] ^ 1);
  assign w610[39] = |(datain[155:152] ^ 15);
  assign w610[40] = |(datain[151:148] ^ 6);
  assign w610[41] = |(datain[147:144] ^ 1);
  assign w610[42] = |(datain[143:140] ^ 14);
  assign w610[43] = |(datain[139:136] ^ 10);
  assign comp[610] = ~(|w610);
  wire [44-1:0] w611;
  assign w611[0] = |(datain[311:308] ^ 4);
  assign w611[1] = |(datain[307:304] ^ 2);
  assign w611[2] = |(datain[303:300] ^ 8);
  assign w611[3] = |(datain[299:296] ^ 11);
  assign w611[4] = |(datain[295:292] ^ 12);
  assign w611[5] = |(datain[291:288] ^ 10);
  assign w611[6] = |(datain[287:284] ^ 12);
  assign w611[7] = |(datain[283:280] ^ 13);
  assign w611[8] = |(datain[279:276] ^ 14);
  assign w611[9] = |(datain[275:272] ^ 5);
  assign w611[10] = |(datain[271:268] ^ 11);
  assign w611[11] = |(datain[267:264] ^ 4);
  assign w611[12] = |(datain[263:260] ^ 4);
  assign w611[13] = |(datain[259:256] ^ 0);
  assign w611[14] = |(datain[255:252] ^ 11);
  assign w611[15] = |(datain[251:248] ^ 2);
  assign w611[16] = |(datain[247:244] ^ 2);
  assign w611[17] = |(datain[243:240] ^ 13);
  assign w611[18] = |(datain[239:236] ^ 11);
  assign w611[19] = |(datain[235:232] ^ 1);
  assign w611[20] = |(datain[231:228] ^ 0);
  assign w611[21] = |(datain[227:224] ^ 3);
  assign w611[22] = |(datain[223:220] ^ 8);
  assign w611[23] = |(datain[219:216] ^ 9);
  assign w611[24] = |(datain[215:212] ^ 2);
  assign w611[25] = |(datain[211:208] ^ 12);
  assign w611[26] = |(datain[207:204] ^ 12);
  assign w611[27] = |(datain[203:200] ^ 13);
  assign w611[28] = |(datain[199:196] ^ 14);
  assign w611[29] = |(datain[195:192] ^ 5);
  assign w611[30] = |(datain[191:188] ^ 11);
  assign w611[31] = |(datain[187:184] ^ 4);
  assign w611[32] = |(datain[183:180] ^ 3);
  assign w611[33] = |(datain[179:176] ^ 14);
  assign w611[34] = |(datain[175:172] ^ 12);
  assign w611[35] = |(datain[171:168] ^ 13);
  assign w611[36] = |(datain[167:164] ^ 14);
  assign w611[37] = |(datain[163:160] ^ 5);
  assign w611[38] = |(datain[159:156] ^ 1);
  assign w611[39] = |(datain[155:152] ^ 15);
  assign w611[40] = |(datain[151:148] ^ 6);
  assign w611[41] = |(datain[147:144] ^ 1);
  assign w611[42] = |(datain[143:140] ^ 14);
  assign w611[43] = |(datain[139:136] ^ 10);
  assign comp[611] = ~(|w611);
  wire [42-1:0] w612;
  assign w612[0] = |(datain[311:308] ^ 8);
  assign w612[1] = |(datain[307:304] ^ 12);
  assign w612[2] = |(datain[303:300] ^ 2);
  assign w612[3] = |(datain[299:296] ^ 11);
  assign w612[4] = |(datain[295:292] ^ 12);
  assign w612[5] = |(datain[291:288] ^ 1);
  assign w612[6] = |(datain[287:284] ^ 3);
  assign w612[7] = |(datain[283:280] ^ 11);
  assign w612[8] = |(datain[279:276] ^ 4);
  assign w612[9] = |(datain[275:272] ^ 4);
  assign w612[10] = |(datain[271:268] ^ 0);
  assign w612[11] = |(datain[267:264] ^ 1);
  assign w612[12] = |(datain[263:260] ^ 7);
  assign w612[13] = |(datain[259:256] ^ 4);
  assign w612[14] = |(datain[255:252] ^ 1);
  assign w612[15] = |(datain[251:248] ^ 6);
  assign w612[16] = |(datain[247:244] ^ 11);
  assign w612[17] = |(datain[243:240] ^ 4);
  assign w612[18] = |(datain[239:236] ^ 4);
  assign w612[19] = |(datain[235:232] ^ 0);
  assign w612[20] = |(datain[231:228] ^ 12);
  assign w612[21] = |(datain[227:224] ^ 13);
  assign w612[22] = |(datain[223:220] ^ 15);
  assign w612[23] = |(datain[219:216] ^ 7);
  assign w612[24] = |(datain[215:212] ^ 11);
  assign w612[25] = |(datain[211:208] ^ 8);
  assign w612[26] = |(datain[207:204] ^ 0);
  assign w612[27] = |(datain[203:200] ^ 0);
  assign w612[28] = |(datain[199:196] ^ 4);
  assign w612[29] = |(datain[195:192] ^ 2);
  assign w612[30] = |(datain[191:188] ^ 3);
  assign w612[31] = |(datain[187:184] ^ 3);
  assign w612[32] = |(datain[183:180] ^ 12);
  assign w612[33] = |(datain[179:176] ^ 9);
  assign w612[34] = |(datain[175:172] ^ 12);
  assign w612[35] = |(datain[171:168] ^ 13);
  assign w612[36] = |(datain[167:164] ^ 15);
  assign w612[37] = |(datain[163:160] ^ 7);
  assign w612[38] = |(datain[159:156] ^ 11);
  assign w612[39] = |(datain[155:152] ^ 4);
  assign w612[40] = |(datain[151:148] ^ 4);
  assign w612[41] = |(datain[147:144] ^ 0);
  assign comp[612] = ~(|w612);
  wire [46-1:0] w613;
  assign w613[0] = |(datain[311:308] ^ 4);
  assign w613[1] = |(datain[307:304] ^ 2);
  assign w613[2] = |(datain[303:300] ^ 3);
  assign w613[3] = |(datain[299:296] ^ 3);
  assign w613[4] = |(datain[295:292] ^ 12);
  assign w613[5] = |(datain[291:288] ^ 9);
  assign w613[6] = |(datain[287:284] ^ 12);
  assign w613[7] = |(datain[283:280] ^ 13);
  assign w613[8] = |(datain[279:276] ^ 11);
  assign w613[9] = |(datain[275:272] ^ 4);
  assign w613[10] = |(datain[271:268] ^ 11);
  assign w613[11] = |(datain[267:264] ^ 4);
  assign w613[12] = |(datain[263:260] ^ 4);
  assign w613[13] = |(datain[259:256] ^ 0);
  assign w613[14] = |(datain[255:252] ^ 8);
  assign w613[15] = |(datain[251:248] ^ 13);
  assign w613[16] = |(datain[247:244] ^ 5);
  assign w613[17] = |(datain[243:240] ^ 4);
  assign w613[18] = |(datain[239:236] ^ 15);
  assign w613[19] = |(datain[235:232] ^ 15);
  assign w613[20] = |(datain[231:228] ^ 11);
  assign w613[21] = |(datain[227:224] ^ 1);
  assign w613[22] = |(datain[223:220] ^ 0);
  assign w613[23] = |(datain[219:216] ^ 3);
  assign w613[24] = |(datain[215:212] ^ 8);
  assign w613[25] = |(datain[211:208] ^ 9);
  assign w613[26] = |(datain[207:204] ^ 2);
  assign w613[27] = |(datain[203:200] ^ 12);
  assign w613[28] = |(datain[199:196] ^ 12);
  assign w613[29] = |(datain[195:192] ^ 13);
  assign w613[30] = |(datain[191:188] ^ 11);
  assign w613[31] = |(datain[187:184] ^ 4);
  assign w613[32] = |(datain[183:180] ^ 11);
  assign w613[33] = |(datain[179:176] ^ 4);
  assign w613[34] = |(datain[175:172] ^ 3);
  assign w613[35] = |(datain[171:168] ^ 14);
  assign w613[36] = |(datain[167:164] ^ 12);
  assign w613[37] = |(datain[163:160] ^ 13);
  assign w613[38] = |(datain[159:156] ^ 11);
  assign w613[39] = |(datain[155:152] ^ 4);
  assign w613[40] = |(datain[151:148] ^ 1);
  assign w613[41] = |(datain[147:144] ^ 15);
  assign w613[42] = |(datain[143:140] ^ 6);
  assign w613[43] = |(datain[139:136] ^ 1);
  assign w613[44] = |(datain[135:132] ^ 14);
  assign w613[45] = |(datain[131:128] ^ 10);
  assign comp[613] = ~(|w613);
  wire [30-1:0] w614;
  assign w614[0] = |(datain[311:308] ^ 10);
  assign w614[1] = |(datain[307:304] ^ 5);
  assign w614[2] = |(datain[303:300] ^ 11);
  assign w614[3] = |(datain[299:296] ^ 8);
  assign w614[4] = |(datain[295:292] ^ 2);
  assign w614[5] = |(datain[291:288] ^ 4);
  assign w614[6] = |(datain[287:284] ^ 0);
  assign w614[7] = |(datain[283:280] ^ 0);
  assign w614[8] = |(datain[279:276] ^ 8);
  assign w614[9] = |(datain[275:272] ^ 14);
  assign w614[10] = |(datain[271:268] ^ 12);
  assign w614[11] = |(datain[267:264] ^ 0);
  assign w614[12] = |(datain[263:260] ^ 3);
  assign w614[13] = |(datain[259:256] ^ 3);
  assign w614[14] = |(datain[255:252] ^ 15);
  assign w614[15] = |(datain[251:248] ^ 15);
  assign w614[16] = |(datain[247:244] ^ 8);
  assign w614[17] = |(datain[243:240] ^ 3);
  assign w614[18] = |(datain[239:236] ^ 14);
  assign w614[19] = |(datain[235:232] ^ 14);
  assign w614[20] = |(datain[231:228] ^ 3);
  assign w614[21] = |(datain[227:224] ^ 10);
  assign w614[22] = |(datain[223:220] ^ 2);
  assign w614[23] = |(datain[219:216] ^ 6);
  assign w614[24] = |(datain[215:212] ^ 8);
  assign w614[25] = |(datain[211:208] ^ 0);
  assign w614[26] = |(datain[207:204] ^ 3);
  assign w614[27] = |(datain[203:200] ^ 13);
  assign w614[28] = |(datain[199:196] ^ 6);
  assign w614[29] = |(datain[195:192] ^ 0);
  assign comp[614] = ~(|w614);
  wire [32-1:0] w615;
  assign w615[0] = |(datain[311:308] ^ 11);
  assign w615[1] = |(datain[307:304] ^ 1);
  assign w615[2] = |(datain[303:300] ^ 9);
  assign w615[3] = |(datain[299:296] ^ 0);
  assign w615[4] = |(datain[295:292] ^ 2);
  assign w615[5] = |(datain[291:288] ^ 11);
  assign w615[6] = |(datain[287:284] ^ 12);
  assign w615[7] = |(datain[283:280] ^ 1);
  assign w615[8] = |(datain[279:276] ^ 3);
  assign w615[9] = |(datain[275:272] ^ 11);
  assign w615[10] = |(datain[271:268] ^ 4);
  assign w615[11] = |(datain[267:264] ^ 4);
  assign w615[12] = |(datain[263:260] ^ 0);
  assign w615[13] = |(datain[259:256] ^ 1);
  assign w615[14] = |(datain[255:252] ^ 7);
  assign w615[15] = |(datain[251:248] ^ 4);
  assign w615[16] = |(datain[247:244] ^ 1);
  assign w615[17] = |(datain[243:240] ^ 6);
  assign w615[18] = |(datain[239:236] ^ 11);
  assign w615[19] = |(datain[235:232] ^ 4);
  assign w615[20] = |(datain[231:228] ^ 4);
  assign w615[21] = |(datain[227:224] ^ 0);
  assign w615[22] = |(datain[223:220] ^ 12);
  assign w615[23] = |(datain[219:216] ^ 13);
  assign w615[24] = |(datain[215:212] ^ 11);
  assign w615[25] = |(datain[211:208] ^ 4);
  assign w615[26] = |(datain[207:204] ^ 11);
  assign w615[27] = |(datain[203:200] ^ 8);
  assign w615[28] = |(datain[199:196] ^ 0);
  assign w615[29] = |(datain[195:192] ^ 0);
  assign w615[30] = |(datain[191:188] ^ 4);
  assign w615[31] = |(datain[187:184] ^ 2);
  assign comp[615] = ~(|w615);
  wire [46-1:0] w616;
  assign w616[0] = |(datain[311:308] ^ 12);
  assign w616[1] = |(datain[307:304] ^ 9);
  assign w616[2] = |(datain[303:300] ^ 3);
  assign w616[3] = |(datain[299:296] ^ 3);
  assign w616[4] = |(datain[295:292] ^ 13);
  assign w616[5] = |(datain[291:288] ^ 2);
  assign w616[6] = |(datain[287:284] ^ 12);
  assign w616[7] = |(datain[283:280] ^ 13);
  assign w616[8] = |(datain[279:276] ^ 2);
  assign w616[9] = |(datain[275:272] ^ 1);
  assign w616[10] = |(datain[271:268] ^ 11);
  assign w616[11] = |(datain[267:264] ^ 4);
  assign w616[12] = |(datain[263:260] ^ 4);
  assign w616[13] = |(datain[259:256] ^ 0);
  assign w616[14] = |(datain[255:252] ^ 8);
  assign w616[15] = |(datain[251:248] ^ 13);
  assign w616[16] = |(datain[247:244] ^ 5);
  assign w616[17] = |(datain[243:240] ^ 4);
  assign w616[18] = |(datain[239:236] ^ 15);
  assign w616[19] = |(datain[235:232] ^ 15);
  assign w616[20] = |(datain[231:228] ^ 11);
  assign w616[21] = |(datain[227:224] ^ 1);
  assign w616[22] = |(datain[223:220] ^ 0);
  assign w616[23] = |(datain[219:216] ^ 3);
  assign w616[24] = |(datain[215:212] ^ 8);
  assign w616[25] = |(datain[211:208] ^ 9);
  assign w616[26] = |(datain[207:204] ^ 2);
  assign w616[27] = |(datain[203:200] ^ 12);
  assign w616[28] = |(datain[199:196] ^ 12);
  assign w616[29] = |(datain[195:192] ^ 13);
  assign w616[30] = |(datain[191:188] ^ 2);
  assign w616[31] = |(datain[187:184] ^ 1);
  assign w616[32] = |(datain[183:180] ^ 11);
  assign w616[33] = |(datain[179:176] ^ 4);
  assign w616[34] = |(datain[175:172] ^ 3);
  assign w616[35] = |(datain[171:168] ^ 14);
  assign w616[36] = |(datain[167:164] ^ 12);
  assign w616[37] = |(datain[163:160] ^ 13);
  assign w616[38] = |(datain[159:156] ^ 2);
  assign w616[39] = |(datain[155:152] ^ 1);
  assign w616[40] = |(datain[151:148] ^ 1);
  assign w616[41] = |(datain[147:144] ^ 15);
  assign w616[42] = |(datain[143:140] ^ 6);
  assign w616[43] = |(datain[139:136] ^ 1);
  assign w616[44] = |(datain[135:132] ^ 14);
  assign w616[45] = |(datain[131:128] ^ 10);
  assign comp[616] = ~(|w616);
  wire [46-1:0] w617;
  assign w617[0] = |(datain[311:308] ^ 10);
  assign w617[1] = |(datain[307:304] ^ 4);
  assign w617[2] = |(datain[303:300] ^ 10);
  assign w617[3] = |(datain[299:296] ^ 5);
  assign w617[4] = |(datain[295:292] ^ 3);
  assign w617[5] = |(datain[291:288] ^ 2);
  assign w617[6] = |(datain[287:284] ^ 12);
  assign w617[7] = |(datain[283:280] ^ 0);
  assign w617[8] = |(datain[279:276] ^ 8);
  assign w617[9] = |(datain[275:272] ^ 14);
  assign w617[10] = |(datain[271:268] ^ 12);
  assign w617[11] = |(datain[267:264] ^ 0);
  assign w617[12] = |(datain[263:260] ^ 11);
  assign w617[13] = |(datain[259:256] ^ 15);
  assign w617[14] = |(datain[255:252] ^ 4);
  assign w617[15] = |(datain[251:248] ^ 0);
  assign w617[16] = |(datain[247:244] ^ 0);
  assign w617[17] = |(datain[243:240] ^ 2);
  assign w617[18] = |(datain[239:236] ^ 8);
  assign w617[19] = |(datain[235:232] ^ 3);
  assign w617[20] = |(datain[231:228] ^ 14);
  assign w617[21] = |(datain[227:224] ^ 14);
  assign w617[22] = |(datain[223:220] ^ 3);
  assign w617[23] = |(datain[219:216] ^ 10);
  assign w617[24] = |(datain[215:212] ^ 2);
  assign w617[25] = |(datain[211:208] ^ 6);
  assign w617[26] = |(datain[207:204] ^ 8);
  assign w617[27] = |(datain[203:200] ^ 0);
  assign w617[28] = |(datain[199:196] ^ 3);
  assign w617[29] = |(datain[195:192] ^ 13);
  assign w617[30] = |(datain[191:188] ^ 6);
  assign w617[31] = |(datain[187:184] ^ 0);
  assign w617[32] = |(datain[183:180] ^ 11);
  assign w617[33] = |(datain[179:176] ^ 1);
  assign w617[34] = |(datain[175:172] ^ 9);
  assign w617[35] = |(datain[171:168] ^ 5);
  assign w617[36] = |(datain[167:164] ^ 15);
  assign w617[37] = |(datain[163:160] ^ 3);
  assign w617[38] = |(datain[159:156] ^ 10);
  assign w617[39] = |(datain[155:152] ^ 4);
  assign w617[40] = |(datain[151:148] ^ 7);
  assign w617[41] = |(datain[147:144] ^ 4);
  assign w617[42] = |(datain[143:140] ^ 1);
  assign w617[43] = |(datain[139:136] ^ 1);
  assign w617[44] = |(datain[135:132] ^ 8);
  assign w617[45] = |(datain[131:128] ^ 14);
  assign comp[617] = ~(|w617);
  wire [42-1:0] w618;
  assign w618[0] = |(datain[311:308] ^ 8);
  assign w618[1] = |(datain[307:304] ^ 11);
  assign w618[2] = |(datain[303:300] ^ 2);
  assign w618[3] = |(datain[299:296] ^ 14);
  assign w618[4] = |(datain[295:292] ^ 0);
  assign w618[5] = |(datain[291:288] ^ 2);
  assign w618[6] = |(datain[287:284] ^ 0);
  assign w618[7] = |(datain[283:280] ^ 1);
  assign w618[8] = |(datain[279:276] ^ 11);
  assign w618[9] = |(datain[275:272] ^ 0);
  assign w618[10] = |(datain[271:268] ^ 0);
  assign w618[11] = |(datain[267:264] ^ 9);
  assign w618[12] = |(datain[263:260] ^ 11);
  assign w618[13] = |(datain[259:256] ^ 9);
  assign w618[14] = |(datain[255:252] ^ 13);
  assign w618[15] = |(datain[251:248] ^ 15);
  assign w618[16] = |(datain[247:244] ^ 0);
  assign w618[17] = |(datain[243:240] ^ 4);
  assign w618[18] = |(datain[239:236] ^ 11);
  assign w618[19] = |(datain[235:232] ^ 14);
  assign w618[20] = |(datain[231:228] ^ 1);
  assign w618[21] = |(datain[227:224] ^ 5);
  assign w618[22] = |(datain[223:220] ^ 0);
  assign w618[23] = |(datain[219:216] ^ 0);
  assign w618[24] = |(datain[215:212] ^ 0);
  assign w618[25] = |(datain[211:208] ^ 1);
  assign w618[26] = |(datain[207:204] ^ 14);
  assign w618[27] = |(datain[203:200] ^ 14);
  assign w618[28] = |(datain[199:196] ^ 3);
  assign w618[29] = |(datain[195:192] ^ 0);
  assign w618[30] = |(datain[191:188] ^ 0);
  assign w618[31] = |(datain[187:184] ^ 4);
  assign w618[32] = |(datain[183:180] ^ 15);
  assign w618[33] = |(datain[179:176] ^ 14);
  assign w618[34] = |(datain[175:172] ^ 12);
  assign w618[35] = |(datain[171:168] ^ 8);
  assign w618[36] = |(datain[167:164] ^ 4);
  assign w618[37] = |(datain[163:160] ^ 6);
  assign w618[38] = |(datain[159:156] ^ 14);
  assign w618[39] = |(datain[155:152] ^ 2);
  assign w618[40] = |(datain[151:148] ^ 15);
  assign w618[41] = |(datain[147:144] ^ 9);
  assign comp[618] = ~(|w618);
  wire [26-1:0] w619;
  assign w619[0] = |(datain[311:308] ^ 8);
  assign w619[1] = |(datain[307:304] ^ 13);
  assign w619[2] = |(datain[303:300] ^ 7);
  assign w619[3] = |(datain[299:296] ^ 12);
  assign w619[4] = |(datain[295:292] ^ 4);
  assign w619[5] = |(datain[291:288] ^ 10);
  assign w619[6] = |(datain[287:284] ^ 15);
  assign w619[7] = |(datain[283:280] ^ 14);
  assign w619[8] = |(datain[279:276] ^ 12);
  assign w619[9] = |(datain[275:272] ^ 2);
  assign w619[10] = |(datain[271:268] ^ 3);
  assign w619[11] = |(datain[267:264] ^ 0);
  assign w619[12] = |(datain[263:260] ^ 1);
  assign w619[13] = |(datain[259:256] ^ 5);
  assign w619[14] = |(datain[255:252] ^ 3);
  assign w619[15] = |(datain[251:248] ^ 0);
  assign w619[16] = |(datain[247:244] ^ 0);
  assign w619[17] = |(datain[243:240] ^ 13);
  assign w619[18] = |(datain[239:236] ^ 4);
  assign w619[19] = |(datain[235:232] ^ 7);
  assign w619[20] = |(datain[231:228] ^ 14);
  assign w619[21] = |(datain[227:224] ^ 2);
  assign w619[22] = |(datain[223:220] ^ 15);
  assign w619[23] = |(datain[219:216] ^ 7);
  assign w619[24] = |(datain[215:212] ^ 12);
  assign w619[25] = |(datain[211:208] ^ 3);
  assign comp[619] = ~(|w619);
  wire [46-1:0] w620;
  assign w620[0] = |(datain[311:308] ^ 3);
  assign w620[1] = |(datain[307:304] ^ 15);
  assign w620[2] = |(datain[303:300] ^ 8);
  assign w620[3] = |(datain[299:296] ^ 13);
  assign w620[4] = |(datain[295:292] ^ 9);
  assign w620[5] = |(datain[291:288] ^ 6);
  assign w620[6] = |(datain[287:284] ^ 8);
  assign w620[7] = |(datain[283:280] ^ 7);
  assign w620[8] = |(datain[279:276] ^ 0);
  assign w620[9] = |(datain[275:272] ^ 0);
  assign w620[10] = |(datain[271:268] ^ 11);
  assign w620[11] = |(datain[267:264] ^ 9);
  assign w620[12] = |(datain[263:260] ^ 0);
  assign w620[13] = |(datain[259:256] ^ 6);
  assign w620[14] = |(datain[255:252] ^ 0);
  assign w620[15] = |(datain[251:248] ^ 0);
  assign w620[16] = |(datain[247:244] ^ 12);
  assign w620[17] = |(datain[243:240] ^ 13);
  assign w620[18] = |(datain[239:236] ^ 2);
  assign w620[19] = |(datain[235:232] ^ 1);
  assign w620[20] = |(datain[231:228] ^ 7);
  assign w620[21] = |(datain[227:224] ^ 2);
  assign w620[22] = |(datain[223:220] ^ 6);
  assign w620[23] = |(datain[219:216] ^ 6);
  assign w620[24] = |(datain[215:212] ^ 11);
  assign w620[25] = |(datain[211:208] ^ 4);
  assign w620[26] = |(datain[207:204] ^ 5);
  assign w620[27] = |(datain[203:200] ^ 10);
  assign w620[28] = |(datain[199:196] ^ 11);
  assign w620[29] = |(datain[195:192] ^ 0);
  assign w620[30] = |(datain[191:188] ^ 4);
  assign w620[31] = |(datain[187:184] ^ 13);
  assign w620[32] = |(datain[183:180] ^ 3);
  assign w620[33] = |(datain[179:176] ^ 9);
  assign w620[34] = |(datain[175:172] ^ 8);
  assign w620[35] = |(datain[171:168] ^ 6);
  assign w620[36] = |(datain[167:164] ^ 8);
  assign w620[37] = |(datain[163:160] ^ 7);
  assign w620[38] = |(datain[159:156] ^ 0);
  assign w620[39] = |(datain[155:152] ^ 0);
  assign w620[40] = |(datain[151:148] ^ 7);
  assign w620[41] = |(datain[147:144] ^ 4);
  assign w620[42] = |(datain[143:140] ^ 0);
  assign w620[43] = |(datain[139:136] ^ 7);
  assign w620[44] = |(datain[135:132] ^ 8);
  assign w620[45] = |(datain[131:128] ^ 0);
  assign comp[620] = ~(|w620);
  wire [44-1:0] w621;
  assign w621[0] = |(datain[311:308] ^ 0);
  assign w621[1] = |(datain[307:304] ^ 5);
  assign w621[2] = |(datain[303:300] ^ 9);
  assign w621[3] = |(datain[299:296] ^ 0);
  assign w621[4] = |(datain[295:292] ^ 11);
  assign w621[5] = |(datain[291:288] ^ 4);
  assign w621[6] = |(datain[287:284] ^ 4);
  assign w621[7] = |(datain[283:280] ^ 0);
  assign w621[8] = |(datain[279:276] ^ 12);
  assign w621[9] = |(datain[275:272] ^ 13);
  assign w621[10] = |(datain[271:268] ^ 2);
  assign w621[11] = |(datain[267:264] ^ 1);
  assign w621[12] = |(datain[263:260] ^ 11);
  assign w621[13] = |(datain[259:256] ^ 4);
  assign w621[14] = |(datain[255:252] ^ 3);
  assign w621[15] = |(datain[251:248] ^ 14);
  assign w621[16] = |(datain[247:244] ^ 12);
  assign w621[17] = |(datain[243:240] ^ 13);
  assign w621[18] = |(datain[239:236] ^ 2);
  assign w621[19] = |(datain[235:232] ^ 1);
  assign w621[20] = |(datain[231:228] ^ 11);
  assign w621[21] = |(datain[227:224] ^ 10);
  assign w621[22] = |(datain[223:220] ^ 14);
  assign w621[23] = |(datain[219:216] ^ 1);
  assign w621[24] = |(datain[215:212] ^ 0);
  assign w621[25] = |(datain[211:208] ^ 0);
  assign w621[26] = |(datain[207:204] ^ 8);
  assign w621[27] = |(datain[203:200] ^ 11);
  assign w621[28] = |(datain[199:196] ^ 0);
  assign w621[29] = |(datain[195:192] ^ 14);
  assign w621[30] = |(datain[191:188] ^ 1);
  assign w621[31] = |(datain[187:184] ^ 12);
  assign w621[32] = |(datain[183:180] ^ 0);
  assign w621[33] = |(datain[179:176] ^ 3);
  assign w621[34] = |(datain[175:172] ^ 15);
  assign w621[35] = |(datain[171:168] ^ 6);
  assign w621[36] = |(datain[167:164] ^ 12);
  assign w621[37] = |(datain[163:160] ^ 1);
  assign w621[38] = |(datain[159:156] ^ 0);
  assign w621[39] = |(datain[155:152] ^ 1);
  assign w621[40] = |(datain[151:148] ^ 7);
  assign w621[41] = |(datain[147:144] ^ 4);
  assign w621[42] = |(datain[143:140] ^ 0);
  assign w621[43] = |(datain[139:136] ^ 5);
  assign comp[621] = ~(|w621);
  wire [40-1:0] w622;
  assign w622[0] = |(datain[311:308] ^ 12);
  assign w622[1] = |(datain[307:304] ^ 0);
  assign w622[2] = |(datain[303:300] ^ 10);
  assign w622[3] = |(datain[299:296] ^ 2);
  assign w622[4] = |(datain[295:292] ^ 0);
  assign w622[5] = |(datain[291:288] ^ 11);
  assign w622[6] = |(datain[287:284] ^ 0);
  assign w622[7] = |(datain[283:280] ^ 0);
  assign w622[8] = |(datain[279:276] ^ 8);
  assign w622[9] = |(datain[275:272] ^ 14);
  assign w622[10] = |(datain[271:268] ^ 13);
  assign w622[11] = |(datain[267:264] ^ 8);
  assign w622[12] = |(datain[263:260] ^ 11);
  assign w622[13] = |(datain[259:256] ^ 0);
  assign w622[14] = |(datain[255:252] ^ 5);
  assign w622[15] = |(datain[251:248] ^ 2);
  assign w622[16] = |(datain[247:244] ^ 10);
  assign w622[17] = |(datain[243:240] ^ 3);
  assign w622[18] = |(datain[239:236] ^ 4);
  assign w622[19] = |(datain[235:232] ^ 12);
  assign w622[20] = |(datain[231:228] ^ 0);
  assign w622[21] = |(datain[227:224] ^ 0);
  assign w622[22] = |(datain[223:220] ^ 8);
  assign w622[23] = |(datain[219:216] ^ 12);
  assign w622[24] = |(datain[215:212] ^ 0);
  assign w622[25] = |(datain[211:208] ^ 14);
  assign w622[26] = |(datain[207:204] ^ 4);
  assign w622[27] = |(datain[203:200] ^ 14);
  assign w622[28] = |(datain[199:196] ^ 0);
  assign w622[29] = |(datain[195:192] ^ 0);
  assign w622[30] = |(datain[191:188] ^ 14);
  assign w622[31] = |(datain[187:184] ^ 10);
  assign w622[32] = |(datain[183:180] ^ 0);
  assign w622[33] = |(datain[179:176] ^ 0);
  assign w622[34] = |(datain[175:172] ^ 0);
  assign w622[35] = |(datain[171:168] ^ 0);
  assign w622[36] = |(datain[167:164] ^ 12);
  assign w622[37] = |(datain[163:160] ^ 0);
  assign w622[38] = |(datain[159:156] ^ 0);
  assign w622[39] = |(datain[155:152] ^ 7);
  assign comp[622] = ~(|w622);
  wire [72-1:0] w623;
  assign w623[0] = |(datain[311:308] ^ 12);
  assign w623[1] = |(datain[307:304] ^ 13);
  assign w623[2] = |(datain[303:300] ^ 2);
  assign w623[3] = |(datain[299:296] ^ 1);
  assign w623[4] = |(datain[295:292] ^ 8);
  assign w623[5] = |(datain[291:288] ^ 12);
  assign w623[6] = |(datain[287:284] ^ 0);
  assign w623[7] = |(datain[283:280] ^ 6);
  assign w623[8] = |(datain[279:276] ^ 6);
  assign w623[9] = |(datain[275:272] ^ 9);
  assign w623[10] = |(datain[271:268] ^ 0);
  assign w623[11] = |(datain[267:264] ^ 0);
  assign w623[12] = |(datain[263:260] ^ 8);
  assign w623[13] = |(datain[259:256] ^ 9);
  assign w623[14] = |(datain[255:252] ^ 1);
  assign w623[15] = |(datain[251:248] ^ 14);
  assign w623[16] = |(datain[247:244] ^ 6);
  assign w623[17] = |(datain[243:240] ^ 7);
  assign w623[18] = |(datain[239:236] ^ 0);
  assign w623[19] = |(datain[235:232] ^ 0);
  assign w623[20] = |(datain[231:228] ^ 11);
  assign w623[21] = |(datain[227:224] ^ 10);
  assign w623[22] = |(datain[223:220] ^ 2);
  assign w623[23] = |(datain[219:216] ^ 0);
  assign w623[24] = |(datain[215:212] ^ 0);
  assign w623[25] = |(datain[211:208] ^ 0);
  assign w623[26] = |(datain[207:204] ^ 8);
  assign w623[27] = |(datain[203:200] ^ 14);
  assign w623[28] = |(datain[199:196] ^ 12);
  assign w623[29] = |(datain[195:192] ^ 2);
  assign w623[30] = |(datain[191:188] ^ 3);
  assign w623[31] = |(datain[187:184] ^ 3);
  assign w623[32] = |(datain[183:180] ^ 15);
  assign w623[33] = |(datain[179:176] ^ 15);
  assign w623[34] = |(datain[175:172] ^ 2);
  assign w623[35] = |(datain[171:168] ^ 6);
  assign w623[36] = |(datain[167:164] ^ 8);
  assign w623[37] = |(datain[163:160] ^ 0);
  assign w623[38] = |(datain[159:156] ^ 3);
  assign w623[39] = |(datain[155:152] ^ 13);
  assign w623[40] = |(datain[151:148] ^ 0);
  assign w623[41] = |(datain[147:144] ^ 6);
  assign w623[42] = |(datain[143:140] ^ 7);
  assign w623[43] = |(datain[139:136] ^ 4);
  assign w623[44] = |(datain[135:132] ^ 0);
  assign w623[45] = |(datain[131:128] ^ 14);
  assign w623[46] = |(datain[127:124] ^ 14);
  assign w623[47] = |(datain[123:120] ^ 8);
  assign w623[48] = |(datain[119:116] ^ 3);
  assign w623[49] = |(datain[115:112] ^ 0);
  assign w623[50] = |(datain[111:108] ^ 0);
  assign w623[51] = |(datain[107:104] ^ 1);
  assign w623[52] = |(datain[103:100] ^ 8);
  assign w623[53] = |(datain[99:96] ^ 14);
  assign w623[54] = |(datain[95:92] ^ 13);
  assign w623[55] = |(datain[91:88] ^ 10);
  assign w623[56] = |(datain[87:84] ^ 11);
  assign w623[57] = |(datain[83:80] ^ 4);
  assign w623[58] = |(datain[79:76] ^ 2);
  assign w623[59] = |(datain[75:72] ^ 5);
  assign w623[60] = |(datain[71:68] ^ 11);
  assign w623[61] = |(datain[67:64] ^ 10);
  assign w623[62] = |(datain[63:60] ^ 5);
  assign w623[63] = |(datain[59:56] ^ 12);
  assign w623[64] = |(datain[55:52] ^ 0);
  assign w623[65] = |(datain[51:48] ^ 0);
  assign w623[66] = |(datain[47:44] ^ 12);
  assign w623[67] = |(datain[43:40] ^ 13);
  assign w623[68] = |(datain[39:36] ^ 2);
  assign w623[69] = |(datain[35:32] ^ 1);
  assign w623[70] = |(datain[31:28] ^ 0);
  assign w623[71] = |(datain[27:24] ^ 14);
  assign comp[623] = ~(|w623);
  wire [42-1:0] w624;
  assign w624[0] = |(datain[311:308] ^ 12);
  assign w624[1] = |(datain[307:304] ^ 13);
  assign w624[2] = |(datain[303:300] ^ 2);
  assign w624[3] = |(datain[299:296] ^ 1);
  assign w624[4] = |(datain[295:292] ^ 3);
  assign w624[5] = |(datain[291:288] ^ 13);
  assign w624[6] = |(datain[287:284] ^ 10);
  assign w624[7] = |(datain[283:280] ^ 1);
  assign w624[8] = |(datain[279:276] ^ 8);
  assign w624[9] = |(datain[275:272] ^ 14);
  assign w624[10] = |(datain[271:268] ^ 7);
  assign w624[11] = |(datain[267:264] ^ 4);
  assign w624[12] = |(datain[263:260] ^ 4);
  assign w624[13] = |(datain[259:256] ^ 4);
  assign w624[14] = |(datain[255:252] ^ 11);
  assign w624[15] = |(datain[251:248] ^ 9);
  assign w624[16] = |(datain[247:244] ^ 2);
  assign w624[17] = |(datain[243:240] ^ 12);
  assign w624[18] = |(datain[239:236] ^ 0);
  assign w624[19] = |(datain[235:232] ^ 1);
  assign w624[20] = |(datain[231:228] ^ 8);
  assign w624[21] = |(datain[227:224] ^ 3);
  assign w624[22] = |(datain[223:220] ^ 2);
  assign w624[23] = |(datain[219:216] ^ 14);
  assign w624[24] = |(datain[215:212] ^ 0);
  assign w624[25] = |(datain[211:208] ^ 2);
  assign w624[26] = |(datain[207:204] ^ 0);
  assign w624[27] = |(datain[203:200] ^ 0);
  assign w624[28] = |(datain[199:196] ^ 1);
  assign w624[29] = |(datain[195:192] ^ 3);
  assign w624[30] = |(datain[191:188] ^ 8);
  assign w624[31] = |(datain[187:184] ^ 12);
  assign w624[32] = |(datain[183:180] ^ 13);
  assign w624[33] = |(datain[179:176] ^ 11);
  assign w624[34] = |(datain[175:172] ^ 4);
  assign w624[35] = |(datain[171:168] ^ 11);
  assign w624[36] = |(datain[167:164] ^ 8);
  assign w624[37] = |(datain[163:160] ^ 14);
  assign w624[38] = |(datain[159:156] ^ 12);
  assign w624[39] = |(datain[155:152] ^ 3);
  assign w624[40] = |(datain[151:148] ^ 2);
  assign w624[41] = |(datain[147:144] ^ 6);
  assign comp[624] = ~(|w624);
  wire [44-1:0] w625;
  assign w625[0] = |(datain[311:308] ^ 5);
  assign w625[1] = |(datain[307:304] ^ 0);
  assign w625[2] = |(datain[303:300] ^ 5);
  assign w625[3] = |(datain[299:296] ^ 3);
  assign w625[4] = |(datain[295:292] ^ 5);
  assign w625[5] = |(datain[291:288] ^ 1);
  assign w625[6] = |(datain[287:284] ^ 14);
  assign w625[7] = |(datain[283:280] ^ 8);
  assign w625[8] = |(datain[279:276] ^ 0);
  assign w625[9] = |(datain[275:272] ^ 1);
  assign w625[10] = |(datain[271:268] ^ 0);
  assign w625[11] = |(datain[267:264] ^ 0);
  assign w625[12] = |(datain[263:260] ^ 7);
  assign w625[13] = |(datain[259:256] ^ 3);
  assign w625[14] = |(datain[255:252] ^ 5);
  assign w625[15] = |(datain[251:248] ^ 13);
  assign w625[16] = |(datain[247:244] ^ 8);
  assign w625[17] = |(datain[243:240] ^ 3);
  assign w625[18] = |(datain[239:236] ^ 14);
  assign w625[19] = |(datain[235:232] ^ 13);
  assign w625[20] = |(datain[231:228] ^ 0);
  assign w625[21] = |(datain[227:224] ^ 8);
  assign w625[22] = |(datain[223:220] ^ 9);
  assign w625[23] = |(datain[219:216] ^ 0);
  assign w625[24] = |(datain[215:212] ^ 15);
  assign w625[25] = |(datain[211:208] ^ 12);
  assign w625[26] = |(datain[207:204] ^ 0);
  assign w625[27] = |(datain[203:200] ^ 14);
  assign w625[28] = |(datain[199:196] ^ 1);
  assign w625[29] = |(datain[195:192] ^ 15);
  assign w625[30] = |(datain[191:188] ^ 11);
  assign w625[31] = |(datain[187:184] ^ 14);
  assign w625[32] = |(datain[183:180] ^ 2);
  assign w625[33] = |(datain[179:176] ^ 8);
  assign w625[34] = |(datain[175:172] ^ 0);
  assign w625[35] = |(datain[171:168] ^ 0);
  assign w625[36] = |(datain[167:164] ^ 0);
  assign w625[37] = |(datain[163:160] ^ 3);
  assign w625[38] = |(datain[159:156] ^ 15);
  assign w625[39] = |(datain[155:152] ^ 5);
  assign w625[40] = |(datain[151:148] ^ 8);
  assign w625[41] = |(datain[147:144] ^ 11);
  assign w625[42] = |(datain[143:140] ^ 15);
  assign w625[43] = |(datain[139:136] ^ 14);
  assign comp[625] = ~(|w625);
  wire [60-1:0] w626;
  assign w626[0] = |(datain[311:308] ^ 8);
  assign w626[1] = |(datain[307:304] ^ 3);
  assign w626[2] = |(datain[303:300] ^ 14);
  assign w626[3] = |(datain[299:296] ^ 13);
  assign w626[4] = |(datain[295:292] ^ 0);
  assign w626[5] = |(datain[291:288] ^ 8);
  assign w626[6] = |(datain[287:284] ^ 15);
  assign w626[7] = |(datain[283:280] ^ 12);
  assign w626[8] = |(datain[279:276] ^ 9);
  assign w626[9] = |(datain[275:272] ^ 0);
  assign w626[10] = |(datain[271:268] ^ 0);
  assign w626[11] = |(datain[267:264] ^ 14);
  assign w626[12] = |(datain[263:260] ^ 11);
  assign w626[13] = |(datain[259:256] ^ 14);
  assign w626[14] = |(datain[255:252] ^ 2);
  assign w626[15] = |(datain[251:248] ^ 8);
  assign w626[16] = |(datain[247:244] ^ 0);
  assign w626[17] = |(datain[243:240] ^ 0);
  assign w626[18] = |(datain[239:236] ^ 1);
  assign w626[19] = |(datain[235:232] ^ 15);
  assign w626[20] = |(datain[231:228] ^ 0);
  assign w626[21] = |(datain[227:224] ^ 3);
  assign w626[22] = |(datain[223:220] ^ 15);
  assign w626[23] = |(datain[219:216] ^ 5);
  assign w626[24] = |(datain[215:212] ^ 8);
  assign w626[25] = |(datain[211:208] ^ 11);
  assign w626[26] = |(datain[207:204] ^ 15);
  assign w626[27] = |(datain[203:200] ^ 14);
  assign w626[28] = |(datain[199:196] ^ 1);
  assign w626[29] = |(datain[195:192] ^ 14);
  assign w626[30] = |(datain[191:188] ^ 11);
  assign w626[31] = |(datain[187:184] ^ 9);
  assign w626[32] = |(datain[183:180] ^ 11);
  assign w626[33] = |(datain[179:176] ^ 8);
  assign w626[34] = |(datain[175:172] ^ 0);
  assign w626[35] = |(datain[171:168] ^ 5);
  assign w626[36] = |(datain[167:164] ^ 0);
  assign w626[37] = |(datain[163:160] ^ 7);
  assign w626[38] = |(datain[159:156] ^ 3);
  assign w626[39] = |(datain[155:152] ^ 14);
  assign w626[40] = |(datain[151:148] ^ 8);
  assign w626[41] = |(datain[147:144] ^ 10);
  assign w626[42] = |(datain[143:140] ^ 6);
  assign w626[43] = |(datain[139:136] ^ 6);
  assign w626[44] = |(datain[135:132] ^ 0);
  assign w626[45] = |(datain[131:128] ^ 8);
  assign w626[46] = |(datain[127:124] ^ 9);
  assign w626[47] = |(datain[123:120] ^ 0);
  assign w626[48] = |(datain[119:116] ^ 10);
  assign w626[49] = |(datain[115:112] ^ 12);
  assign w626[50] = |(datain[111:108] ^ 3);
  assign w626[51] = |(datain[107:104] ^ 2);
  assign w626[52] = |(datain[103:100] ^ 12);
  assign w626[53] = |(datain[99:96] ^ 4);
  assign w626[54] = |(datain[95:92] ^ 10);
  assign w626[55] = |(datain[91:88] ^ 10);
  assign w626[56] = |(datain[87:84] ^ 14);
  assign w626[57] = |(datain[83:80] ^ 2);
  assign w626[58] = |(datain[79:76] ^ 15);
  assign w626[59] = |(datain[75:72] ^ 10);
  assign comp[626] = ~(|w626);
  wire [58-1:0] w627;
  assign w627[0] = |(datain[311:308] ^ 14);
  assign w627[1] = |(datain[307:304] ^ 13);
  assign w627[2] = |(datain[303:300] ^ 0);
  assign w627[3] = |(datain[299:296] ^ 8);
  assign w627[4] = |(datain[295:292] ^ 9);
  assign w627[5] = |(datain[291:288] ^ 0);
  assign w627[6] = |(datain[287:284] ^ 15);
  assign w627[7] = |(datain[283:280] ^ 12);
  assign w627[8] = |(datain[279:276] ^ 0);
  assign w627[9] = |(datain[275:272] ^ 14);
  assign w627[10] = |(datain[271:268] ^ 1);
  assign w627[11] = |(datain[267:264] ^ 15);
  assign w627[12] = |(datain[263:260] ^ 11);
  assign w627[13] = |(datain[259:256] ^ 14);
  assign w627[14] = |(datain[255:252] ^ 2);
  assign w627[15] = |(datain[251:248] ^ 8);
  assign w627[16] = |(datain[247:244] ^ 0);
  assign w627[17] = |(datain[243:240] ^ 0);
  assign w627[18] = |(datain[239:236] ^ 0);
  assign w627[19] = |(datain[235:232] ^ 3);
  assign w627[20] = |(datain[231:228] ^ 15);
  assign w627[21] = |(datain[227:224] ^ 5);
  assign w627[22] = |(datain[223:220] ^ 8);
  assign w627[23] = |(datain[219:216] ^ 11);
  assign w627[24] = |(datain[215:212] ^ 15);
  assign w627[25] = |(datain[211:208] ^ 14);
  assign w627[26] = |(datain[207:204] ^ 1);
  assign w627[27] = |(datain[203:200] ^ 14);
  assign w627[28] = |(datain[199:196] ^ 0);
  assign w627[29] = |(datain[195:192] ^ 7);
  assign w627[30] = |(datain[191:188] ^ 11);
  assign w627[31] = |(datain[187:184] ^ 9);
  assign w627[32] = |(datain[183:180] ^ 15);
  assign w627[33] = |(datain[179:176] ^ 1);
  assign w627[34] = |(datain[175:172] ^ 0);
  assign w627[35] = |(datain[171:168] ^ 5);
  assign w627[36] = |(datain[167:164] ^ 3);
  assign w627[37] = |(datain[163:160] ^ 14);
  assign w627[38] = |(datain[159:156] ^ 8);
  assign w627[39] = |(datain[155:152] ^ 10);
  assign w627[40] = |(datain[151:148] ^ 9);
  assign w627[41] = |(datain[147:144] ^ 14);
  assign w627[42] = |(datain[143:140] ^ 0);
  assign w627[43] = |(datain[139:136] ^ 8);
  assign w627[44] = |(datain[135:132] ^ 0);
  assign w627[45] = |(datain[131:128] ^ 0);
  assign w627[46] = |(datain[127:124] ^ 10);
  assign w627[47] = |(datain[123:120] ^ 12);
  assign w627[48] = |(datain[119:116] ^ 3);
  assign w627[49] = |(datain[115:112] ^ 2);
  assign w627[50] = |(datain[111:108] ^ 12);
  assign w627[51] = |(datain[107:104] ^ 3);
  assign w627[52] = |(datain[103:100] ^ 10);
  assign w627[53] = |(datain[99:96] ^ 10);
  assign w627[54] = |(datain[95:92] ^ 14);
  assign w627[55] = |(datain[91:88] ^ 2);
  assign w627[56] = |(datain[87:84] ^ 15);
  assign w627[57] = |(datain[83:80] ^ 10);
  assign comp[627] = ~(|w627);
  wire [44-1:0] w628;
  assign w628[0] = |(datain[311:308] ^ 0);
  assign w628[1] = |(datain[307:304] ^ 14);
  assign w628[2] = |(datain[303:300] ^ 0);
  assign w628[3] = |(datain[299:296] ^ 14);
  assign w628[4] = |(datain[295:292] ^ 10);
  assign w628[5] = |(datain[291:288] ^ 15);
  assign w628[6] = |(datain[287:284] ^ 11);
  assign w628[7] = |(datain[283:280] ^ 0);
  assign w628[8] = |(datain[279:276] ^ 2);
  assign w628[9] = |(datain[275:272] ^ 7);
  assign w628[10] = |(datain[271:268] ^ 11);
  assign w628[11] = |(datain[267:264] ^ 3);
  assign w628[12] = |(datain[263:260] ^ 1);
  assign w628[13] = |(datain[259:256] ^ 4);
  assign w628[14] = |(datain[255:252] ^ 8);
  assign w628[15] = |(datain[251:248] ^ 14);
  assign w628[16] = |(datain[247:244] ^ 12);
  assign w628[17] = |(datain[243:240] ^ 0);
  assign w628[18] = |(datain[239:236] ^ 6);
  assign w628[19] = |(datain[235:232] ^ 0);
  assign w628[20] = |(datain[231:228] ^ 10);
  assign w628[21] = |(datain[227:224] ^ 7);
  assign w628[22] = |(datain[223:220] ^ 6);
  assign w628[23] = |(datain[219:216] ^ 1);
  assign w628[24] = |(datain[215:212] ^ 11);
  assign w628[25] = |(datain[211:208] ^ 1);
  assign w628[26] = |(datain[207:204] ^ 7);
  assign w628[27] = |(datain[203:200] ^ 0);
  assign w628[28] = |(datain[199:196] ^ 15);
  assign w628[29] = |(datain[195:192] ^ 3);
  assign w628[30] = |(datain[191:188] ^ 10);
  assign w628[31] = |(datain[187:184] ^ 4);
  assign w628[32] = |(datain[183:180] ^ 8);
  assign w628[33] = |(datain[179:176] ^ 14);
  assign w628[34] = |(datain[175:172] ^ 13);
  assign w628[35] = |(datain[171:168] ^ 9);
  assign w628[36] = |(datain[167:164] ^ 7);
  assign w628[37] = |(datain[163:160] ^ 4);
  assign w628[38] = |(datain[159:156] ^ 0);
  assign w628[39] = |(datain[155:152] ^ 8);
  assign w628[40] = |(datain[151:148] ^ 5);
  assign w628[41] = |(datain[147:144] ^ 0);
  assign w628[42] = |(datain[143:140] ^ 8);
  assign w628[43] = |(datain[139:136] ^ 7);
  assign comp[628] = ~(|w628);
  wire [42-1:0] w629;
  assign w629[0] = |(datain[311:308] ^ 0);
  assign w629[1] = |(datain[307:304] ^ 6);
  assign w629[2] = |(datain[303:300] ^ 8);
  assign w629[3] = |(datain[299:296] ^ 0);
  assign w629[4] = |(datain[295:292] ^ 15);
  assign w629[5] = |(datain[291:288] ^ 4);
  assign w629[6] = |(datain[287:284] ^ 4);
  assign w629[7] = |(datain[283:280] ^ 11);
  assign w629[8] = |(datain[279:276] ^ 7);
  assign w629[9] = |(datain[275:272] ^ 5);
  assign w629[10] = |(datain[271:268] ^ 3);
  assign w629[11] = |(datain[267:264] ^ 13);
  assign w629[12] = |(datain[263:260] ^ 11);
  assign w629[13] = |(datain[259:256] ^ 8);
  assign w629[14] = |(datain[255:252] ^ 0);
  assign w629[15] = |(datain[251:248] ^ 2);
  assign w629[16] = |(datain[247:244] ^ 3);
  assign w629[17] = |(datain[243:240] ^ 13);
  assign w629[18] = |(datain[239:236] ^ 12);
  assign w629[19] = |(datain[235:232] ^ 13);
  assign w629[20] = |(datain[231:228] ^ 12);
  assign w629[21] = |(datain[227:224] ^ 5);
  assign w629[22] = |(datain[223:220] ^ 7);
  assign w629[23] = |(datain[219:216] ^ 2);
  assign w629[24] = |(datain[215:212] ^ 3);
  assign w629[25] = |(datain[211:208] ^ 6);
  assign w629[26] = |(datain[207:204] ^ 9);
  assign w629[27] = |(datain[203:200] ^ 3);
  assign w629[28] = |(datain[199:196] ^ 3);
  assign w629[29] = |(datain[195:192] ^ 3);
  assign w629[30] = |(datain[191:188] ^ 15);
  assign w629[31] = |(datain[187:184] ^ 15);
  assign w629[32] = |(datain[183:180] ^ 11);
  assign w629[33] = |(datain[179:176] ^ 5);
  assign w629[34] = |(datain[175:172] ^ 8);
  assign w629[35] = |(datain[171:168] ^ 12);
  assign w629[36] = |(datain[167:164] ^ 8);
  assign w629[37] = |(datain[163:160] ^ 14);
  assign w629[38] = |(datain[159:156] ^ 13);
  assign w629[39] = |(datain[155:152] ^ 9);
  assign w629[40] = |(datain[151:148] ^ 1);
  assign w629[41] = |(datain[147:144] ^ 14);
  assign comp[629] = ~(|w629);
  wire [46-1:0] w630;
  assign w630[0] = |(datain[311:308] ^ 0);
  assign w630[1] = |(datain[307:304] ^ 14);
  assign w630[2] = |(datain[303:300] ^ 5);
  assign w630[3] = |(datain[299:296] ^ 6);
  assign w630[4] = |(datain[295:292] ^ 0);
  assign w630[5] = |(datain[291:288] ^ 14);
  assign w630[6] = |(datain[287:284] ^ 11);
  assign w630[7] = |(datain[283:280] ^ 0);
  assign w630[8] = |(datain[279:276] ^ 2);
  assign w630[9] = |(datain[275:272] ^ 14);
  assign w630[10] = |(datain[271:268] ^ 5);
  assign w630[11] = |(datain[267:264] ^ 0);
  assign w630[12] = |(datain[263:260] ^ 8);
  assign w630[13] = |(datain[259:256] ^ 14);
  assign w630[14] = |(datain[255:252] ^ 12);
  assign w630[15] = |(datain[251:248] ^ 0);
  assign w630[16] = |(datain[247:244] ^ 3);
  assign w630[17] = |(datain[243:240] ^ 3);
  assign w630[18] = |(datain[239:236] ^ 15);
  assign w630[19] = |(datain[235:232] ^ 15);
  assign w630[20] = |(datain[231:228] ^ 11);
  assign w630[21] = |(datain[227:224] ^ 1);
  assign w630[22] = |(datain[223:220] ^ 7);
  assign w630[23] = |(datain[219:216] ^ 8);
  assign w630[24] = |(datain[215:212] ^ 15);
  assign w630[25] = |(datain[211:208] ^ 3);
  assign w630[26] = |(datain[207:204] ^ 10);
  assign w630[27] = |(datain[203:200] ^ 4);
  assign w630[28] = |(datain[199:196] ^ 6);
  assign w630[29] = |(datain[195:192] ^ 10);
  assign w630[30] = |(datain[191:188] ^ 1);
  assign w630[31] = |(datain[187:184] ^ 2);
  assign w630[32] = |(datain[183:180] ^ 12);
  assign w630[33] = |(datain[179:176] ^ 11);
  assign w630[34] = |(datain[175:172] ^ 5);
  assign w630[35] = |(datain[171:168] ^ 6);
  assign w630[36] = |(datain[167:164] ^ 11);
  assign w630[37] = |(datain[163:160] ^ 14);
  assign w630[38] = |(datain[159:156] ^ 8);
  assign w630[39] = |(datain[155:152] ^ 4);
  assign w630[40] = |(datain[151:148] ^ 0);
  assign w630[41] = |(datain[147:144] ^ 0);
  assign w630[42] = |(datain[143:140] ^ 8);
  assign w630[43] = |(datain[139:136] ^ 14);
  assign w630[44] = |(datain[135:132] ^ 13);
  assign w630[45] = |(datain[131:128] ^ 9);
  assign comp[630] = ~(|w630);
  wire [74-1:0] w631;
  assign w631[0] = |(datain[311:308] ^ 9);
  assign w631[1] = |(datain[307:304] ^ 14);
  assign w631[2] = |(datain[303:300] ^ 5);
  assign w631[3] = |(datain[299:296] ^ 8);
  assign w631[4] = |(datain[295:292] ^ 0);
  assign w631[5] = |(datain[291:288] ^ 2);
  assign w631[6] = |(datain[287:284] ^ 8);
  assign w631[7] = |(datain[283:280] ^ 9);
  assign w631[8] = |(datain[279:276] ^ 0);
  assign w631[9] = |(datain[275:272] ^ 7);
  assign w631[10] = |(datain[271:268] ^ 5);
  assign w631[11] = |(datain[267:264] ^ 11);
  assign w631[12] = |(datain[263:260] ^ 11);
  assign w631[13] = |(datain[259:256] ^ 4);
  assign w631[14] = |(datain[255:252] ^ 4);
  assign w631[15] = |(datain[251:248] ^ 0);
  assign w631[16] = |(datain[247:244] ^ 11);
  assign w631[17] = |(datain[243:240] ^ 9);
  assign w631[18] = |(datain[239:236] ^ 5);
  assign w631[19] = |(datain[235:232] ^ 14);
  assign w631[20] = |(datain[231:228] ^ 0);
  assign w631[21] = |(datain[227:224] ^ 1);
  assign w631[22] = |(datain[223:220] ^ 8);
  assign w631[23] = |(datain[219:216] ^ 13);
  assign w631[24] = |(datain[215:212] ^ 9);
  assign w631[25] = |(datain[211:208] ^ 6);
  assign w631[26] = |(datain[207:204] ^ 0);
  assign w631[27] = |(datain[203:200] ^ 5);
  assign w631[28] = |(datain[199:196] ^ 0);
  assign w631[29] = |(datain[195:192] ^ 1);
  assign w631[30] = |(datain[191:188] ^ 12);
  assign w631[31] = |(datain[187:184] ^ 13);
  assign w631[32] = |(datain[183:180] ^ 2);
  assign w631[33] = |(datain[179:176] ^ 1);
  assign w631[34] = |(datain[175:172] ^ 11);
  assign w631[35] = |(datain[171:168] ^ 8);
  assign w631[36] = |(datain[167:164] ^ 0);
  assign w631[37] = |(datain[163:160] ^ 0);
  assign w631[38] = |(datain[159:156] ^ 4);
  assign w631[39] = |(datain[155:152] ^ 2);
  assign w631[40] = |(datain[151:148] ^ 3);
  assign w631[41] = |(datain[147:144] ^ 3);
  assign w631[42] = |(datain[143:140] ^ 12);
  assign w631[43] = |(datain[139:136] ^ 9);
  assign w631[44] = |(datain[135:132] ^ 3);
  assign w631[45] = |(datain[131:128] ^ 3);
  assign w631[46] = |(datain[127:124] ^ 13);
  assign w631[47] = |(datain[123:120] ^ 2);
  assign w631[48] = |(datain[119:116] ^ 12);
  assign w631[49] = |(datain[115:112] ^ 13);
  assign w631[50] = |(datain[111:108] ^ 2);
  assign w631[51] = |(datain[107:104] ^ 1);
  assign w631[52] = |(datain[103:100] ^ 11);
  assign w631[53] = |(datain[99:96] ^ 4);
  assign w631[54] = |(datain[95:92] ^ 4);
  assign w631[55] = |(datain[91:88] ^ 0);
  assign w631[56] = |(datain[87:84] ^ 11);
  assign w631[57] = |(datain[83:80] ^ 9);
  assign w631[58] = |(datain[79:76] ^ 0);
  assign w631[59] = |(datain[75:72] ^ 1);
  assign w631[60] = |(datain[71:68] ^ 0);
  assign w631[61] = |(datain[67:64] ^ 0);
  assign w631[62] = |(datain[63:60] ^ 8);
  assign w631[63] = |(datain[59:56] ^ 13);
  assign w631[64] = |(datain[55:52] ^ 9);
  assign w631[65] = |(datain[51:48] ^ 6);
  assign w631[66] = |(datain[47:44] ^ 5);
  assign w631[67] = |(datain[43:40] ^ 7);
  assign w631[68] = |(datain[39:36] ^ 0);
  assign w631[69] = |(datain[35:32] ^ 2);
  assign w631[70] = |(datain[31:28] ^ 12);
  assign w631[71] = |(datain[27:24] ^ 13);
  assign w631[72] = |(datain[23:20] ^ 2);
  assign w631[73] = |(datain[19:16] ^ 1);
  assign comp[631] = ~(|w631);
  wire [74-1:0] w632;
  assign w632[0] = |(datain[311:308] ^ 0);
  assign w632[1] = |(datain[307:304] ^ 2);
  assign w632[2] = |(datain[303:300] ^ 3);
  assign w632[3] = |(datain[299:296] ^ 13);
  assign w632[4] = |(datain[295:292] ^ 11);
  assign w632[5] = |(datain[291:288] ^ 10);
  assign w632[6] = |(datain[287:284] ^ 9);
  assign w632[7] = |(datain[283:280] ^ 14);
  assign w632[8] = |(datain[279:276] ^ 0);
  assign w632[9] = |(datain[275:272] ^ 0);
  assign w632[10] = |(datain[271:268] ^ 12);
  assign w632[11] = |(datain[267:264] ^ 13);
  assign w632[12] = |(datain[263:260] ^ 2);
  assign w632[13] = |(datain[259:256] ^ 1);
  assign w632[14] = |(datain[255:252] ^ 9);
  assign w632[15] = |(datain[251:248] ^ 3);
  assign w632[16] = |(datain[247:244] ^ 11);
  assign w632[17] = |(datain[243:240] ^ 8);
  assign w632[18] = |(datain[239:236] ^ 0);
  assign w632[19] = |(datain[235:232] ^ 0);
  assign w632[20] = |(datain[231:228] ^ 5);
  assign w632[21] = |(datain[227:224] ^ 7);
  assign w632[22] = |(datain[223:220] ^ 12);
  assign w632[23] = |(datain[219:216] ^ 13);
  assign w632[24] = |(datain[215:212] ^ 2);
  assign w632[25] = |(datain[211:208] ^ 1);
  assign w632[26] = |(datain[207:204] ^ 5);
  assign w632[27] = |(datain[203:200] ^ 2);
  assign w632[28] = |(datain[199:196] ^ 5);
  assign w632[29] = |(datain[195:192] ^ 1);
  assign w632[30] = |(datain[191:188] ^ 11);
  assign w632[31] = |(datain[187:184] ^ 4);
  assign w632[32] = |(datain[183:180] ^ 4);
  assign w632[33] = |(datain[179:176] ^ 0);
  assign w632[34] = |(datain[175:172] ^ 11);
  assign w632[35] = |(datain[171:168] ^ 9);
  assign w632[36] = |(datain[167:164] ^ 7);
  assign w632[37] = |(datain[163:160] ^ 3);
  assign w632[38] = |(datain[159:156] ^ 0);
  assign w632[39] = |(datain[155:152] ^ 1);
  assign w632[40] = |(datain[151:148] ^ 11);
  assign w632[41] = |(datain[147:144] ^ 10);
  assign w632[42] = |(datain[143:140] ^ 0);
  assign w632[43] = |(datain[139:136] ^ 0);
  assign w632[44] = |(datain[135:132] ^ 0);
  assign w632[45] = |(datain[131:128] ^ 1);
  assign w632[46] = |(datain[127:124] ^ 12);
  assign w632[47] = |(datain[123:120] ^ 13);
  assign w632[48] = |(datain[119:116] ^ 2);
  assign w632[49] = |(datain[115:112] ^ 1);
  assign w632[50] = |(datain[111:108] ^ 11);
  assign w632[51] = |(datain[107:104] ^ 8);
  assign w632[52] = |(datain[103:100] ^ 0);
  assign w632[53] = |(datain[99:96] ^ 1);
  assign w632[54] = |(datain[95:92] ^ 5);
  assign w632[55] = |(datain[91:88] ^ 7);
  assign w632[56] = |(datain[87:84] ^ 5);
  assign w632[57] = |(datain[83:80] ^ 9);
  assign w632[58] = |(datain[79:76] ^ 5);
  assign w632[59] = |(datain[75:72] ^ 10);
  assign w632[60] = |(datain[71:68] ^ 12);
  assign w632[61] = |(datain[67:64] ^ 13);
  assign w632[62] = |(datain[63:60] ^ 2);
  assign w632[63] = |(datain[59:56] ^ 1);
  assign w632[64] = |(datain[55:52] ^ 11);
  assign w632[65] = |(datain[51:48] ^ 4);
  assign w632[66] = |(datain[47:44] ^ 3);
  assign w632[67] = |(datain[43:40] ^ 14);
  assign w632[68] = |(datain[39:36] ^ 12);
  assign w632[69] = |(datain[35:32] ^ 13);
  assign w632[70] = |(datain[31:28] ^ 2);
  assign w632[71] = |(datain[27:24] ^ 1);
  assign w632[72] = |(datain[23:20] ^ 12);
  assign w632[73] = |(datain[19:16] ^ 3);
  assign comp[632] = ~(|w632);
  wire [54-1:0] w633;
  assign w633[0] = |(datain[311:308] ^ 14);
  assign w633[1] = |(datain[307:304] ^ 8);
  assign w633[2] = |(datain[303:300] ^ 0);
  assign w633[3] = |(datain[299:296] ^ 0);
  assign w633[4] = |(datain[295:292] ^ 0);
  assign w633[5] = |(datain[291:288] ^ 0);
  assign w633[6] = |(datain[287:284] ^ 5);
  assign w633[7] = |(datain[283:280] ^ 13);
  assign w633[8] = |(datain[279:276] ^ 5);
  assign w633[9] = |(datain[275:272] ^ 1);
  assign w633[10] = |(datain[271:268] ^ 5);
  assign w633[11] = |(datain[267:264] ^ 0);
  assign w633[12] = |(datain[263:260] ^ 2);
  assign w633[13] = |(datain[259:256] ^ 14);
  assign w633[14] = |(datain[255:252] ^ 8);
  assign w633[15] = |(datain[251:248] ^ 11);
  assign w633[16] = |(datain[247:244] ^ 4);
  assign w633[17] = |(datain[243:240] ^ 6);
  assign w633[18] = |(datain[239:236] ^ 15);
  assign w633[19] = |(datain[235:232] ^ 10);
  assign w633[20] = |(datain[231:228] ^ 8);
  assign w633[21] = |(datain[227:224] ^ 11);
  assign w633[22] = |(datain[223:220] ^ 15);
  assign w633[23] = |(datain[219:216] ^ 5);
  assign w633[24] = |(datain[215:212] ^ 8);
  assign w633[25] = |(datain[211:208] ^ 3);
  assign w633[26] = |(datain[207:204] ^ 12);
  assign w633[27] = |(datain[203:200] ^ 6);
  assign w633[28] = |(datain[199:196] ^ 1);
  assign w633[29] = |(datain[195:192] ^ 8);
  assign w633[30] = |(datain[191:188] ^ 11);
  assign w633[31] = |(datain[187:184] ^ 9);
  assign w633[32] = |(datain[183:180] ^ 4);
  assign w633[33] = |(datain[179:176] ^ 1);
  assign w633[34] = |(datain[175:172] ^ 0);
  assign w633[35] = |(datain[171:168] ^ 8);
  assign w633[36] = |(datain[167:164] ^ 2);
  assign w633[37] = |(datain[163:160] ^ 14);
  assign w633[38] = |(datain[159:156] ^ 3);
  assign w633[39] = |(datain[155:152] ^ 0);
  assign w633[40] = |(datain[151:148] ^ 0);
  assign w633[41] = |(datain[147:144] ^ 4);
  assign w633[42] = |(datain[143:140] ^ 2);
  assign w633[43] = |(datain[139:136] ^ 14);
  assign w633[44] = |(datain[135:132] ^ 0);
  assign w633[45] = |(datain[131:128] ^ 0);
  assign w633[46] = |(datain[127:124] ^ 2);
  assign w633[47] = |(datain[123:120] ^ 4);
  assign w633[48] = |(datain[119:116] ^ 4);
  assign w633[49] = |(datain[115:112] ^ 6);
  assign w633[50] = |(datain[111:108] ^ 14);
  assign w633[51] = |(datain[107:104] ^ 2);
  assign w633[52] = |(datain[103:100] ^ 15);
  assign w633[53] = |(datain[99:96] ^ 7);
  assign comp[633] = ~(|w633);
  wire [44-1:0] w634;
  assign w634[0] = |(datain[311:308] ^ 4);
  assign w634[1] = |(datain[307:304] ^ 11);
  assign w634[2] = |(datain[303:300] ^ 7);
  assign w634[3] = |(datain[299:296] ^ 4);
  assign w634[4] = |(datain[295:292] ^ 3);
  assign w634[5] = |(datain[291:288] ^ 15);
  assign w634[6] = |(datain[287:284] ^ 3);
  assign w634[7] = |(datain[283:280] ^ 13);
  assign w634[8] = |(datain[279:276] ^ 15);
  assign w634[9] = |(datain[275:272] ^ 15);
  assign w634[10] = |(datain[271:268] ^ 3);
  assign w634[11] = |(datain[267:264] ^ 5);
  assign w634[12] = |(datain[263:260] ^ 7);
  assign w634[13] = |(datain[259:256] ^ 4);
  assign w634[14] = |(datain[255:252] ^ 0);
  assign w634[15] = |(datain[251:248] ^ 15);
  assign w634[16] = |(datain[247:244] ^ 8);
  assign w634[17] = |(datain[243:240] ^ 0);
  assign w634[18] = |(datain[239:236] ^ 15);
  assign w634[19] = |(datain[235:232] ^ 12);
  assign w634[20] = |(datain[231:228] ^ 4);
  assign w634[21] = |(datain[227:224] ^ 1);
  assign w634[22] = |(datain[223:220] ^ 7);
  assign w634[23] = |(datain[219:216] ^ 4);
  assign w634[24] = |(datain[215:212] ^ 0);
  assign w634[25] = |(datain[211:208] ^ 15);
  assign w634[26] = |(datain[207:204] ^ 8);
  assign w634[27] = |(datain[203:200] ^ 0);
  assign w634[28] = |(datain[199:196] ^ 15);
  assign w634[29] = |(datain[195:192] ^ 12);
  assign w634[30] = |(datain[191:188] ^ 1);
  assign w634[31] = |(datain[187:184] ^ 3);
  assign w634[32] = |(datain[183:180] ^ 7);
  assign w634[33] = |(datain[179:176] ^ 4);
  assign w634[34] = |(datain[175:172] ^ 0);
  assign w634[35] = |(datain[171:168] ^ 10);
  assign w634[36] = |(datain[167:164] ^ 2);
  assign w634[37] = |(datain[163:160] ^ 14);
  assign w634[38] = |(datain[159:156] ^ 15);
  assign w634[39] = |(datain[155:152] ^ 15);
  assign w634[40] = |(datain[151:148] ^ 2);
  assign w634[41] = |(datain[147:144] ^ 14);
  assign w634[42] = |(datain[143:140] ^ 14);
  assign w634[43] = |(datain[139:136] ^ 12);
  assign comp[634] = ~(|w634);
  wire [76-1:0] w635;
  assign w635[0] = |(datain[311:308] ^ 12);
  assign w635[1] = |(datain[307:304] ^ 13);
  assign w635[2] = |(datain[303:300] ^ 2);
  assign w635[3] = |(datain[299:296] ^ 1);
  assign w635[4] = |(datain[295:292] ^ 12);
  assign w635[5] = |(datain[291:288] ^ 3);
  assign w635[6] = |(datain[287:284] ^ 11);
  assign w635[7] = |(datain[283:280] ^ 0);
  assign w635[8] = |(datain[279:276] ^ 0);
  assign w635[9] = |(datain[275:272] ^ 2);
  assign w635[10] = |(datain[271:268] ^ 11);
  assign w635[11] = |(datain[267:264] ^ 10);
  assign w635[12] = |(datain[263:260] ^ 9);
  assign w635[13] = |(datain[259:256] ^ 14);
  assign w635[14] = |(datain[255:252] ^ 0);
  assign w635[15] = |(datain[251:248] ^ 0);
  assign w635[16] = |(datain[247:244] ^ 14);
  assign w635[17] = |(datain[243:240] ^ 8);
  assign w635[18] = |(datain[239:236] ^ 14);
  assign w635[19] = |(datain[235:232] ^ 12);
  assign w635[20] = |(datain[231:228] ^ 15);
  assign w635[21] = |(datain[227:224] ^ 15);
  assign w635[22] = |(datain[223:220] ^ 7);
  assign w635[23] = |(datain[219:216] ^ 2);
  assign w635[24] = |(datain[215:212] ^ 2);
  assign w635[25] = |(datain[211:208] ^ 10);
  assign w635[26] = |(datain[207:204] ^ 9);
  assign w635[27] = |(datain[203:200] ^ 3);
  assign w635[28] = |(datain[199:196] ^ 11);
  assign w635[29] = |(datain[195:192] ^ 0);
  assign w635[30] = |(datain[191:188] ^ 0);
  assign w635[31] = |(datain[187:184] ^ 0);
  assign w635[32] = |(datain[183:180] ^ 14);
  assign w635[33] = |(datain[179:176] ^ 8);
  assign w635[34] = |(datain[175:172] ^ 14);
  assign w635[35] = |(datain[171:168] ^ 11);
  assign w635[36] = |(datain[167:164] ^ 15);
  assign w635[37] = |(datain[163:160] ^ 15);
  assign w635[38] = |(datain[159:156] ^ 5);
  assign w635[39] = |(datain[155:152] ^ 1);
  assign w635[40] = |(datain[151:148] ^ 5);
  assign w635[41] = |(datain[147:144] ^ 2);
  assign w635[42] = |(datain[143:140] ^ 11);
  assign w635[43] = |(datain[139:136] ^ 4);
  assign w635[44] = |(datain[135:132] ^ 4);
  assign w635[45] = |(datain[131:128] ^ 0);
  assign w635[46] = |(datain[127:124] ^ 11);
  assign w635[47] = |(datain[123:120] ^ 9);
  assign w635[48] = |(datain[119:116] ^ 14);
  assign w635[49] = |(datain[115:112] ^ 8);
  assign w635[50] = |(datain[111:108] ^ 0);
  assign w635[51] = |(datain[107:104] ^ 0);
  assign w635[52] = |(datain[103:100] ^ 11);
  assign w635[53] = |(datain[99:96] ^ 10);
  assign w635[54] = |(datain[95:92] ^ 0);
  assign w635[55] = |(datain[91:88] ^ 0);
  assign w635[56] = |(datain[87:84] ^ 0);
  assign w635[57] = |(datain[83:80] ^ 1);
  assign w635[58] = |(datain[79:76] ^ 12);
  assign w635[59] = |(datain[75:72] ^ 13);
  assign w635[60] = |(datain[71:68] ^ 2);
  assign w635[61] = |(datain[67:64] ^ 1);
  assign w635[62] = |(datain[63:60] ^ 11);
  assign w635[63] = |(datain[59:56] ^ 0);
  assign w635[64] = |(datain[55:52] ^ 0);
  assign w635[65] = |(datain[51:48] ^ 1);
  assign w635[66] = |(datain[47:44] ^ 5);
  assign w635[67] = |(datain[43:40] ^ 10);
  assign w635[68] = |(datain[39:36] ^ 5);
  assign w635[69] = |(datain[35:32] ^ 9);
  assign w635[70] = |(datain[31:28] ^ 14);
  assign w635[71] = |(datain[27:24] ^ 8);
  assign w635[72] = |(datain[23:20] ^ 13);
  assign w635[73] = |(datain[19:16] ^ 8);
  assign w635[74] = |(datain[15:12] ^ 15);
  assign w635[75] = |(datain[11:8] ^ 15);
  assign comp[635] = ~(|w635);
  wire [76-1:0] w636;
  assign w636[0] = |(datain[311:308] ^ 0);
  assign w636[1] = |(datain[307:304] ^ 7);
  assign w636[2] = |(datain[303:300] ^ 0);
  assign w636[3] = |(datain[299:296] ^ 1);
  assign w636[4] = |(datain[295:292] ^ 11);
  assign w636[5] = |(datain[291:288] ^ 8);
  assign w636[6] = |(datain[287:284] ^ 0);
  assign w636[7] = |(datain[283:280] ^ 2);
  assign w636[8] = |(datain[279:276] ^ 4);
  assign w636[9] = |(datain[275:272] ^ 2);
  assign w636[10] = |(datain[271:268] ^ 3);
  assign w636[11] = |(datain[267:264] ^ 3);
  assign w636[12] = |(datain[263:260] ^ 12);
  assign w636[13] = |(datain[259:256] ^ 9);
  assign w636[14] = |(datain[255:252] ^ 3);
  assign w636[15] = |(datain[251:248] ^ 3);
  assign w636[16] = |(datain[247:244] ^ 13);
  assign w636[17] = |(datain[243:240] ^ 2);
  assign w636[18] = |(datain[239:236] ^ 12);
  assign w636[19] = |(datain[235:232] ^ 13);
  assign w636[20] = |(datain[231:228] ^ 2);
  assign w636[21] = |(datain[227:224] ^ 1);
  assign w636[22] = |(datain[223:220] ^ 11);
  assign w636[23] = |(datain[219:216] ^ 10);
  assign w636[24] = |(datain[215:212] ^ 0);
  assign w636[25] = |(datain[211:208] ^ 12);
  assign w636[26] = |(datain[207:204] ^ 0);
  assign w636[27] = |(datain[203:200] ^ 1);
  assign w636[28] = |(datain[199:196] ^ 11);
  assign w636[29] = |(datain[195:192] ^ 9);
  assign w636[30] = |(datain[191:188] ^ 1);
  assign w636[31] = |(datain[187:184] ^ 15);
  assign w636[32] = |(datain[183:180] ^ 0);
  assign w636[33] = |(datain[179:176] ^ 0);
  assign w636[34] = |(datain[175:172] ^ 11);
  assign w636[35] = |(datain[171:168] ^ 4);
  assign w636[36] = |(datain[167:164] ^ 4);
  assign w636[37] = |(datain[163:160] ^ 0);
  assign w636[38] = |(datain[159:156] ^ 12);
  assign w636[39] = |(datain[155:152] ^ 13);
  assign w636[40] = |(datain[151:148] ^ 2);
  assign w636[41] = |(datain[147:144] ^ 1);
  assign w636[42] = |(datain[143:140] ^ 14);
  assign w636[43] = |(datain[139:136] ^ 9);
  assign w636[44] = |(datain[135:132] ^ 5);
  assign w636[45] = |(datain[131:128] ^ 9);
  assign w636[46] = |(datain[127:124] ^ 0);
  assign w636[47] = |(datain[123:120] ^ 0);
  assign w636[48] = |(datain[119:116] ^ 5);
  assign w636[49] = |(datain[115:112] ^ 14);
  assign w636[50] = |(datain[111:108] ^ 1);
  assign w636[51] = |(datain[107:104] ^ 15);
  assign w636[52] = |(datain[103:100] ^ 0);
  assign w636[53] = |(datain[99:96] ^ 14);
  assign w636[54] = |(datain[95:92] ^ 0);
  assign w636[55] = |(datain[91:88] ^ 7);
  assign w636[56] = |(datain[87:84] ^ 11);
  assign w636[57] = |(datain[83:80] ^ 15);
  assign w636[58] = |(datain[79:76] ^ 2);
  assign w636[59] = |(datain[75:72] ^ 11);
  assign w636[60] = |(datain[71:68] ^ 0);
  assign w636[61] = |(datain[67:64] ^ 1);
  assign w636[62] = |(datain[63:60] ^ 11);
  assign w636[63] = |(datain[59:56] ^ 9);
  assign w636[64] = |(datain[55:52] ^ 4);
  assign w636[65] = |(datain[51:48] ^ 0);
  assign w636[66] = |(datain[47:44] ^ 0);
  assign w636[67] = |(datain[43:40] ^ 0);
  assign w636[68] = |(datain[39:36] ^ 15);
  assign w636[69] = |(datain[35:32] ^ 3);
  assign w636[70] = |(datain[31:28] ^ 10);
  assign w636[71] = |(datain[27:24] ^ 4);
  assign w636[72] = |(datain[23:20] ^ 0);
  assign w636[73] = |(datain[19:16] ^ 14);
  assign w636[74] = |(datain[15:12] ^ 1);
  assign w636[75] = |(datain[11:8] ^ 15);
  assign comp[636] = ~(|w636);
  wire [70-1:0] w637;
  assign w637[0] = |(datain[311:308] ^ 9);
  assign w637[1] = |(datain[307:304] ^ 6);
  assign w637[2] = |(datain[303:300] ^ 2);
  assign w637[3] = |(datain[299:296] ^ 9);
  assign w637[4] = |(datain[295:292] ^ 0);
  assign w637[5] = |(datain[291:288] ^ 3);
  assign w637[6] = |(datain[287:284] ^ 12);
  assign w637[7] = |(datain[283:280] ^ 13);
  assign w637[8] = |(datain[279:276] ^ 2);
  assign w637[9] = |(datain[275:272] ^ 1);
  assign w637[10] = |(datain[271:268] ^ 11);
  assign w637[11] = |(datain[267:264] ^ 9);
  assign w637[12] = |(datain[263:260] ^ 15);
  assign w637[13] = |(datain[259:256] ^ 15);
  assign w637[14] = |(datain[255:252] ^ 1);
  assign w637[15] = |(datain[251:248] ^ 15);
  assign w637[16] = |(datain[247:244] ^ 14);
  assign w637[17] = |(datain[243:240] ^ 2);
  assign w637[18] = |(datain[239:236] ^ 15);
  assign w637[19] = |(datain[235:232] ^ 14);
  assign w637[20] = |(datain[231:228] ^ 14);
  assign w637[21] = |(datain[227:224] ^ 10);
  assign w637[22] = |(datain[223:220] ^ 0);
  assign w637[23] = |(datain[219:216] ^ 0);
  assign w637[24] = |(datain[215:212] ^ 0);
  assign w637[25] = |(datain[211:208] ^ 0);
  assign w637[26] = |(datain[207:204] ^ 15);
  assign w637[27] = |(datain[203:200] ^ 15);
  assign w637[28] = |(datain[199:196] ^ 15);
  assign w637[29] = |(datain[195:192] ^ 15);
  assign w637[30] = |(datain[191:188] ^ 11);
  assign w637[31] = |(datain[187:184] ^ 4);
  assign w637[32] = |(datain[183:180] ^ 1);
  assign w637[33] = |(datain[179:176] ^ 10);
  assign w637[34] = |(datain[175:172] ^ 12);
  assign w637[35] = |(datain[171:168] ^ 13);
  assign w637[36] = |(datain[167:164] ^ 2);
  assign w637[37] = |(datain[163:160] ^ 1);
  assign w637[38] = |(datain[159:156] ^ 12);
  assign w637[39] = |(datain[155:152] ^ 3);
  assign w637[40] = |(datain[151:148] ^ 11);
  assign w637[41] = |(datain[147:144] ^ 4);
  assign w637[42] = |(datain[143:140] ^ 5);
  assign w637[43] = |(datain[139:136] ^ 7);
  assign w637[44] = |(datain[135:132] ^ 12);
  assign w637[45] = |(datain[131:128] ^ 13);
  assign w637[46] = |(datain[127:124] ^ 2);
  assign w637[47] = |(datain[123:120] ^ 1);
  assign w637[48] = |(datain[119:116] ^ 12);
  assign w637[49] = |(datain[115:112] ^ 3);
  assign w637[50] = |(datain[111:108] ^ 11);
  assign w637[51] = |(datain[107:104] ^ 4);
  assign w637[52] = |(datain[103:100] ^ 4);
  assign w637[53] = |(datain[99:96] ^ 3);
  assign w637[54] = |(datain[95:92] ^ 12);
  assign w637[55] = |(datain[91:88] ^ 13);
  assign w637[56] = |(datain[87:84] ^ 2);
  assign w637[57] = |(datain[83:80] ^ 1);
  assign w637[58] = |(datain[79:76] ^ 12);
  assign w637[59] = |(datain[75:72] ^ 3);
  assign w637[60] = |(datain[71:68] ^ 11);
  assign w637[61] = |(datain[67:64] ^ 4);
  assign w637[62] = |(datain[63:60] ^ 4);
  assign w637[63] = |(datain[59:56] ^ 2);
  assign w637[64] = |(datain[55:52] ^ 12);
  assign w637[65] = |(datain[51:48] ^ 13);
  assign w637[66] = |(datain[47:44] ^ 2);
  assign w637[67] = |(datain[43:40] ^ 1);
  assign w637[68] = |(datain[39:36] ^ 12);
  assign w637[69] = |(datain[35:32] ^ 3);
  assign comp[637] = ~(|w637);
  wire [28-1:0] w638;
  assign w638[0] = |(datain[311:308] ^ 0);
  assign w638[1] = |(datain[307:304] ^ 3);
  assign w638[2] = |(datain[303:300] ^ 0);
  assign w638[3] = |(datain[299:296] ^ 0);
  assign w638[4] = |(datain[295:292] ^ 11);
  assign w638[5] = |(datain[291:288] ^ 10);
  assign w638[6] = |(datain[287:284] ^ 7);
  assign w638[7] = |(datain[283:280] ^ 7);
  assign w638[8] = |(datain[279:276] ^ 0);
  assign w638[9] = |(datain[275:272] ^ 2);
  assign w638[10] = |(datain[271:268] ^ 8);
  assign w638[11] = |(datain[267:264] ^ 11);
  assign w638[12] = |(datain[263:260] ^ 15);
  assign w638[13] = |(datain[259:256] ^ 2);
  assign w638[14] = |(datain[255:252] ^ 12);
  assign w638[15] = |(datain[251:248] ^ 13);
  assign w638[16] = |(datain[247:244] ^ 2);
  assign w638[17] = |(datain[243:240] ^ 1);
  assign w638[18] = |(datain[239:236] ^ 8);
  assign w638[19] = |(datain[235:232] ^ 0);
  assign w638[20] = |(datain[231:228] ^ 3);
  assign w638[21] = |(datain[227:224] ^ 12);
  assign w638[22] = |(datain[223:220] ^ 4);
  assign w638[23] = |(datain[219:216] ^ 13);
  assign w638[24] = |(datain[215:212] ^ 7);
  assign w638[25] = |(datain[211:208] ^ 4);
  assign w638[26] = |(datain[207:204] ^ 3);
  assign w638[27] = |(datain[203:200] ^ 1);
  assign comp[638] = ~(|w638);
  wire [42-1:0] w639;
  assign w639[0] = |(datain[311:308] ^ 8);
  assign w639[1] = |(datain[307:304] ^ 3);
  assign w639[2] = |(datain[303:300] ^ 14);
  assign w639[3] = |(datain[299:296] ^ 14);
  assign w639[4] = |(datain[295:292] ^ 3);
  assign w639[5] = |(datain[291:288] ^ 10);
  assign w639[6] = |(datain[287:284] ^ 2);
  assign w639[7] = |(datain[283:280] ^ 6);
  assign w639[8] = |(datain[279:276] ^ 8);
  assign w639[9] = |(datain[275:272] ^ 0);
  assign w639[10] = |(datain[271:268] ^ 3);
  assign w639[11] = |(datain[267:264] ^ 13);
  assign w639[12] = |(datain[263:260] ^ 6);
  assign w639[13] = |(datain[259:256] ^ 0);
  assign w639[14] = |(datain[255:252] ^ 11);
  assign w639[15] = |(datain[251:248] ^ 1);
  assign w639[16] = |(datain[247:244] ^ 9);
  assign w639[17] = |(datain[243:240] ^ 5);
  assign w639[18] = |(datain[239:236] ^ 15);
  assign w639[19] = |(datain[235:232] ^ 3);
  assign w639[20] = |(datain[231:228] ^ 10);
  assign w639[21] = |(datain[227:224] ^ 4);
  assign w639[22] = |(datain[223:220] ^ 7);
  assign w639[23] = |(datain[219:216] ^ 4);
  assign w639[24] = |(datain[215:212] ^ 1);
  assign w639[25] = |(datain[211:208] ^ 1);
  assign w639[26] = |(datain[207:204] ^ 8);
  assign w639[27] = |(datain[203:200] ^ 14);
  assign w639[28] = |(datain[199:196] ^ 13);
  assign w639[29] = |(datain[195:192] ^ 8);
  assign w639[30] = |(datain[191:188] ^ 11);
  assign w639[31] = |(datain[187:184] ^ 14);
  assign w639[32] = |(datain[183:180] ^ 8);
  assign w639[33] = |(datain[179:176] ^ 4);
  assign w639[34] = |(datain[175:172] ^ 0);
  assign w639[35] = |(datain[171:168] ^ 0);
  assign w639[36] = |(datain[167:164] ^ 10);
  assign w639[37] = |(datain[163:160] ^ 5);
  assign w639[38] = |(datain[159:156] ^ 10);
  assign w639[39] = |(datain[155:152] ^ 5);
  assign w639[40] = |(datain[151:148] ^ 12);
  assign w639[41] = |(datain[147:144] ^ 7);
  assign comp[639] = ~(|w639);
  wire [74-1:0] w640;
  assign w640[0] = |(datain[311:308] ^ 11);
  assign w640[1] = |(datain[307:304] ^ 9);
  assign w640[2] = |(datain[303:300] ^ 0);
  assign w640[3] = |(datain[299:296] ^ 3);
  assign w640[4] = |(datain[295:292] ^ 0);
  assign w640[5] = |(datain[291:288] ^ 0);
  assign w640[6] = |(datain[287:284] ^ 5);
  assign w640[7] = |(datain[283:280] ^ 14);
  assign w640[8] = |(datain[279:276] ^ 5);
  assign w640[9] = |(datain[275:272] ^ 15);
  assign w640[10] = |(datain[271:268] ^ 5);
  assign w640[11] = |(datain[267:264] ^ 7);
  assign w640[12] = |(datain[263:260] ^ 5);
  assign w640[13] = |(datain[259:256] ^ 6);
  assign w640[14] = |(datain[255:252] ^ 11);
  assign w640[15] = |(datain[251:248] ^ 10);
  assign w640[16] = |(datain[247:244] ^ 2);
  assign w640[17] = |(datain[243:240] ^ 0);
  assign w640[18] = |(datain[239:236] ^ 0);
  assign w640[19] = |(datain[235:232] ^ 13);
  assign w640[20] = |(datain[231:228] ^ 0);
  assign w640[21] = |(datain[227:224] ^ 3);
  assign w640[22] = |(datain[223:220] ^ 13);
  assign w640[23] = |(datain[219:216] ^ 6);
  assign w640[24] = |(datain[215:212] ^ 1);
  assign w640[25] = |(datain[211:208] ^ 14);
  assign w640[26] = |(datain[207:204] ^ 8);
  assign w640[27] = |(datain[203:200] ^ 14);
  assign w640[28] = |(datain[199:196] ^ 13);
  assign w640[29] = |(datain[195:192] ^ 15);
  assign w640[30] = |(datain[191:188] ^ 12);
  assign w640[31] = |(datain[187:184] ^ 13);
  assign w640[32] = |(datain[183:180] ^ 2);
  assign w640[33] = |(datain[179:176] ^ 1);
  assign w640[34] = |(datain[175:172] ^ 1);
  assign w640[35] = |(datain[171:168] ^ 15);
  assign w640[36] = |(datain[167:164] ^ 11);
  assign w640[37] = |(datain[163:160] ^ 4);
  assign w640[38] = |(datain[159:156] ^ 4);
  assign w640[39] = |(datain[155:152] ^ 2);
  assign w640[40] = |(datain[151:148] ^ 11);
  assign w640[41] = |(datain[147:144] ^ 0);
  assign w640[42] = |(datain[143:140] ^ 0);
  assign w640[43] = |(datain[139:136] ^ 2);
  assign w640[44] = |(datain[135:132] ^ 11);
  assign w640[45] = |(datain[131:128] ^ 9);
  assign w640[46] = |(datain[127:124] ^ 0);
  assign w640[47] = |(datain[123:120] ^ 0);
  assign w640[48] = |(datain[119:116] ^ 0);
  assign w640[49] = |(datain[115:112] ^ 0);
  assign w640[50] = |(datain[111:108] ^ 11);
  assign w640[51] = |(datain[107:104] ^ 10);
  assign w640[52] = |(datain[103:100] ^ 0);
  assign w640[53] = |(datain[99:96] ^ 0);
  assign w640[54] = |(datain[95:92] ^ 0);
  assign w640[55] = |(datain[91:88] ^ 0);
  assign w640[56] = |(datain[87:84] ^ 12);
  assign w640[57] = |(datain[83:80] ^ 13);
  assign w640[58] = |(datain[79:76] ^ 2);
  assign w640[59] = |(datain[75:72] ^ 1);
  assign w640[60] = |(datain[71:68] ^ 0);
  assign w640[61] = |(datain[67:64] ^ 6);
  assign w640[62] = |(datain[63:60] ^ 1);
  assign w640[63] = |(datain[59:56] ^ 15);
  assign w640[64] = |(datain[55:52] ^ 11);
  assign w640[65] = |(datain[51:48] ^ 4);
  assign w640[66] = |(datain[47:44] ^ 4);
  assign w640[67] = |(datain[43:40] ^ 0);
  assign w640[68] = |(datain[39:36] ^ 11);
  assign w640[69] = |(datain[35:32] ^ 9);
  assign w640[70] = |(datain[31:28] ^ 0);
  assign w640[71] = |(datain[27:24] ^ 0);
  assign w640[72] = |(datain[23:20] ^ 0);
  assign w640[73] = |(datain[19:16] ^ 14);
  assign comp[640] = ~(|w640);
  wire [28-1:0] w641;
  assign w641[0] = |(datain[311:308] ^ 8);
  assign w641[1] = |(datain[307:304] ^ 11);
  assign w641[2] = |(datain[303:300] ^ 4);
  assign w641[3] = |(datain[299:296] ^ 7);
  assign w641[4] = |(datain[295:292] ^ 0);
  assign w641[5] = |(datain[291:288] ^ 2);
  assign w641[6] = |(datain[287:284] ^ 8);
  assign w641[7] = |(datain[283:280] ^ 12);
  assign w641[8] = |(datain[279:276] ^ 4);
  assign w641[9] = |(datain[275:272] ^ 7);
  assign w641[10] = |(datain[271:268] ^ 0);
  assign w641[11] = |(datain[267:264] ^ 2);
  assign w641[12] = |(datain[263:260] ^ 2);
  assign w641[13] = |(datain[259:256] ^ 6);
  assign w641[14] = |(datain[255:252] ^ 10);
  assign w641[15] = |(datain[251:248] ^ 3);
  assign w641[16] = |(datain[247:244] ^ 1);
  assign w641[17] = |(datain[243:240] ^ 7);
  assign w641[18] = |(datain[239:236] ^ 0);
  assign w641[19] = |(datain[235:232] ^ 0);
  assign w641[20] = |(datain[231:228] ^ 8);
  assign w641[21] = |(datain[227:224] ^ 12);
  assign w641[22] = |(datain[223:220] ^ 0);
  assign w641[23] = |(datain[219:216] ^ 6);
  assign w641[24] = |(datain[215:212] ^ 1);
  assign w641[25] = |(datain[211:208] ^ 5);
  assign w641[26] = |(datain[207:204] ^ 0);
  assign w641[27] = |(datain[203:200] ^ 4);
  assign comp[641] = ~(|w641);
  wire [32-1:0] w642;
  assign w642[0] = |(datain[311:308] ^ 11);
  assign w642[1] = |(datain[307:304] ^ 0);
  assign w642[2] = |(datain[303:300] ^ 0);
  assign w642[3] = |(datain[299:296] ^ 0);
  assign w642[4] = |(datain[295:292] ^ 8);
  assign w642[5] = |(datain[291:288] ^ 11);
  assign w642[6] = |(datain[287:284] ^ 13);
  assign w642[7] = |(datain[283:280] ^ 10);
  assign w642[8] = |(datain[279:276] ^ 11);
  assign w642[9] = |(datain[275:272] ^ 5);
  assign w642[10] = |(datain[271:268] ^ 0);
  assign w642[11] = |(datain[267:264] ^ 1);
  assign w642[12] = |(datain[263:260] ^ 4);
  assign w642[13] = |(datain[259:256] ^ 3);
  assign w642[14] = |(datain[255:252] ^ 3);
  assign w642[15] = |(datain[251:248] ^ 10);
  assign w642[16] = |(datain[247:244] ^ 0);
  assign w642[17] = |(datain[243:240] ^ 7);
  assign w642[18] = |(datain[239:236] ^ 7);
  assign w642[19] = |(datain[235:232] ^ 5);
  assign w642[20] = |(datain[231:228] ^ 15);
  assign w642[21] = |(datain[227:224] ^ 11);
  assign w642[22] = |(datain[223:220] ^ 4);
  assign w642[23] = |(datain[219:216] ^ 11);
  assign w642[24] = |(datain[215:212] ^ 4);
  assign w642[25] = |(datain[211:208] ^ 11);
  assign w642[26] = |(datain[207:204] ^ 8);
  assign w642[27] = |(datain[203:200] ^ 1);
  assign w642[28] = |(datain[199:196] ^ 2);
  assign w642[29] = |(datain[195:192] ^ 7);
  assign w642[30] = |(datain[191:188] ^ 5);
  assign w642[31] = |(datain[187:184] ^ 15);
  assign comp[642] = ~(|w642);
  wire [44-1:0] w643;
  assign w643[0] = |(datain[311:308] ^ 11);
  assign w643[1] = |(datain[307:304] ^ 8);
  assign w643[2] = |(datain[303:300] ^ 0);
  assign w643[3] = |(datain[299:296] ^ 1);
  assign w643[4] = |(datain[295:292] ^ 15);
  assign w643[5] = |(datain[291:288] ^ 10);
  assign w643[6] = |(datain[287:284] ^ 11);
  assign w643[7] = |(datain[283:280] ^ 10);
  assign w643[8] = |(datain[279:276] ^ 4);
  assign w643[9] = |(datain[275:272] ^ 5);
  assign w643[10] = |(datain[271:268] ^ 5);
  assign w643[11] = |(datain[267:264] ^ 9);
  assign w643[12] = |(datain[263:260] ^ 12);
  assign w643[13] = |(datain[259:256] ^ 13);
  assign w643[14] = |(datain[255:252] ^ 1);
  assign w643[15] = |(datain[251:248] ^ 6);
  assign w643[16] = |(datain[247:244] ^ 14);
  assign w643[17] = |(datain[243:240] ^ 8);
  assign w643[18] = |(datain[239:236] ^ 0);
  assign w643[19] = |(datain[235:232] ^ 0);
  assign w643[20] = |(datain[231:228] ^ 0);
  assign w643[21] = |(datain[227:224] ^ 0);
  assign w643[22] = |(datain[223:220] ^ 5);
  assign w643[23] = |(datain[219:216] ^ 13);
  assign w643[24] = |(datain[215:212] ^ 8);
  assign w643[25] = |(datain[211:208] ^ 1);
  assign w643[26] = |(datain[207:204] ^ 14);
  assign w643[27] = |(datain[203:200] ^ 13);
  assign w643[28] = |(datain[199:196] ^ 0);
  assign w643[29] = |(datain[195:192] ^ 13);
  assign w643[30] = |(datain[191:188] ^ 0);
  assign w643[31] = |(datain[187:184] ^ 1);
  assign w643[32] = |(datain[183:180] ^ 8);
  assign w643[33] = |(datain[179:176] ^ 11);
  assign w643[34] = |(datain[175:172] ^ 12);
  assign w643[35] = |(datain[171:168] ^ 5);
  assign w643[36] = |(datain[167:164] ^ 0);
  assign w643[37] = |(datain[163:160] ^ 5);
  assign w643[38] = |(datain[159:156] ^ 1);
  assign w643[39] = |(datain[155:152] ^ 10);
  assign w643[40] = |(datain[151:148] ^ 0);
  assign w643[41] = |(datain[147:144] ^ 1);
  assign w643[42] = |(datain[143:140] ^ 5);
  assign w643[43] = |(datain[139:136] ^ 0);
  assign comp[643] = ~(|w643);
  wire [38-1:0] w644;
  assign w644[0] = |(datain[311:308] ^ 2);
  assign w644[1] = |(datain[307:304] ^ 6);
  assign w644[2] = |(datain[303:300] ^ 0);
  assign w644[3] = |(datain[299:296] ^ 0);
  assign w644[4] = |(datain[295:292] ^ 15);
  assign w644[5] = |(datain[291:288] ^ 12);
  assign w644[6] = |(datain[287:284] ^ 8);
  assign w644[7] = |(datain[283:280] ^ 10);
  assign w644[8] = |(datain[279:276] ^ 2);
  assign w644[9] = |(datain[275:272] ^ 6);
  assign w644[10] = |(datain[271:268] ^ 0);
  assign w644[11] = |(datain[267:264] ^ 14);
  assign w644[12] = |(datain[263:260] ^ 0);
  assign w644[13] = |(datain[259:256] ^ 0);
  assign w644[14] = |(datain[255:252] ^ 11);
  assign w644[15] = |(datain[251:248] ^ 9);
  assign w644[16] = |(datain[247:244] ^ 6);
  assign w644[17] = |(datain[243:240] ^ 7);
  assign w644[18] = |(datain[239:236] ^ 0);
  assign w644[19] = |(datain[235:232] ^ 2);
  assign w644[20] = |(datain[231:228] ^ 8);
  assign w644[21] = |(datain[227:224] ^ 10);
  assign w644[22] = |(datain[223:220] ^ 0);
  assign w644[23] = |(datain[219:216] ^ 4);
  assign w644[24] = |(datain[215:212] ^ 3);
  assign w644[25] = |(datain[211:208] ^ 2);
  assign w644[26] = |(datain[207:204] ^ 12);
  assign w644[27] = |(datain[203:200] ^ 4);
  assign w644[28] = |(datain[199:196] ^ 8);
  assign w644[29] = |(datain[195:192] ^ 8);
  assign w644[30] = |(datain[191:188] ^ 0);
  assign w644[31] = |(datain[187:184] ^ 4);
  assign w644[32] = |(datain[183:180] ^ 4);
  assign w644[33] = |(datain[179:176] ^ 6);
  assign w644[34] = |(datain[175:172] ^ 14);
  assign w644[35] = |(datain[171:168] ^ 2);
  assign w644[36] = |(datain[167:164] ^ 15);
  assign w644[37] = |(datain[163:160] ^ 7);
  assign comp[644] = ~(|w644);
  wire [40-1:0] w645;
  assign w645[0] = |(datain[311:308] ^ 11);
  assign w645[1] = |(datain[307:304] ^ 4);
  assign w645[2] = |(datain[303:300] ^ 4);
  assign w645[3] = |(datain[299:296] ^ 0);
  assign w645[4] = |(datain[295:292] ^ 11);
  assign w645[5] = |(datain[291:288] ^ 1);
  assign w645[6] = |(datain[287:284] ^ 9);
  assign w645[7] = |(datain[283:280] ^ 3);
  assign w645[8] = |(datain[279:276] ^ 11);
  assign w645[9] = |(datain[275:272] ^ 10);
  assign w645[10] = |(datain[271:268] ^ 0);
  assign w645[11] = |(datain[267:264] ^ 0);
  assign w645[12] = |(datain[263:260] ^ 0);
  assign w645[13] = |(datain[259:256] ^ 1);
  assign w645[14] = |(datain[255:252] ^ 12);
  assign w645[15] = |(datain[251:248] ^ 13);
  assign w645[16] = |(datain[247:244] ^ 2);
  assign w645[17] = |(datain[243:240] ^ 1);
  assign w645[18] = |(datain[239:236] ^ 11);
  assign w645[19] = |(datain[235:232] ^ 4);
  assign w645[20] = |(datain[231:228] ^ 3);
  assign w645[21] = |(datain[227:224] ^ 14);
  assign w645[22] = |(datain[223:220] ^ 12);
  assign w645[23] = |(datain[219:216] ^ 13);
  assign w645[24] = |(datain[215:212] ^ 2);
  assign w645[25] = |(datain[211:208] ^ 1);
  assign w645[26] = |(datain[207:204] ^ 11);
  assign w645[27] = |(datain[203:200] ^ 4);
  assign w645[28] = |(datain[199:196] ^ 4);
  assign w645[29] = |(datain[195:192] ^ 15);
  assign w645[30] = |(datain[191:188] ^ 12);
  assign w645[31] = |(datain[187:184] ^ 13);
  assign w645[32] = |(datain[183:180] ^ 2);
  assign w645[33] = |(datain[179:176] ^ 1);
  assign w645[34] = |(datain[175:172] ^ 7);
  assign w645[35] = |(datain[171:168] ^ 3);
  assign w645[36] = |(datain[167:164] ^ 13);
  assign w645[37] = |(datain[163:160] ^ 3);
  assign w645[38] = |(datain[159:156] ^ 12);
  assign w645[39] = |(datain[155:152] ^ 3);
  assign comp[645] = ~(|w645);
  wire [44-1:0] w646;
  assign w646[0] = |(datain[311:308] ^ 0);
  assign w646[1] = |(datain[307:304] ^ 1);
  assign w646[2] = |(datain[303:300] ^ 11);
  assign w646[3] = |(datain[299:296] ^ 4);
  assign w646[4] = |(datain[295:292] ^ 4);
  assign w646[5] = |(datain[291:288] ^ 0);
  assign w646[6] = |(datain[287:284] ^ 11);
  assign w646[7] = |(datain[283:280] ^ 9);
  assign w646[8] = |(datain[279:276] ^ 4);
  assign w646[9] = |(datain[275:272] ^ 9);
  assign w646[10] = |(datain[271:268] ^ 0);
  assign w646[11] = |(datain[267:264] ^ 5);
  assign w646[12] = |(datain[263:260] ^ 8);
  assign w646[13] = |(datain[259:256] ^ 13);
  assign w646[14] = |(datain[255:252] ^ 9);
  assign w646[15] = |(datain[251:248] ^ 6);
  assign w646[16] = |(datain[247:244] ^ 0);
  assign w646[17] = |(datain[243:240] ^ 0);
  assign w646[18] = |(datain[239:236] ^ 0);
  assign w646[19] = |(datain[235:232] ^ 1);
  assign w646[20] = |(datain[231:228] ^ 12);
  assign w646[21] = |(datain[227:224] ^ 13);
  assign w646[22] = |(datain[223:220] ^ 2);
  assign w646[23] = |(datain[219:216] ^ 1);
  assign w646[24] = |(datain[215:212] ^ 11);
  assign w646[25] = |(datain[211:208] ^ 8);
  assign w646[26] = |(datain[207:204] ^ 0);
  assign w646[27] = |(datain[203:200] ^ 0);
  assign w646[28] = |(datain[199:196] ^ 4);
  assign w646[29] = |(datain[195:192] ^ 2);
  assign w646[30] = |(datain[191:188] ^ 3);
  assign w646[31] = |(datain[187:184] ^ 3);
  assign w646[32] = |(datain[183:180] ^ 12);
  assign w646[33] = |(datain[179:176] ^ 9);
  assign w646[34] = |(datain[175:172] ^ 9);
  assign w646[35] = |(datain[171:168] ^ 9);
  assign w646[36] = |(datain[167:164] ^ 12);
  assign w646[37] = |(datain[163:160] ^ 13);
  assign w646[38] = |(datain[159:156] ^ 2);
  assign w646[39] = |(datain[155:152] ^ 1);
  assign w646[40] = |(datain[151:148] ^ 11);
  assign w646[41] = |(datain[147:144] ^ 4);
  assign w646[42] = |(datain[143:140] ^ 4);
  assign w646[43] = |(datain[139:136] ^ 0);
  assign comp[646] = ~(|w646);
  wire [40-1:0] w647;
  assign w647[0] = |(datain[311:308] ^ 11);
  assign w647[1] = |(datain[307:304] ^ 10);
  assign w647[2] = |(datain[303:300] ^ 6);
  assign w647[3] = |(datain[299:296] ^ 13);
  assign w647[4] = |(datain[295:292] ^ 5);
  assign w647[5] = |(datain[291:288] ^ 4);
  assign w647[6] = |(datain[287:284] ^ 0);
  assign w647[7] = |(datain[283:280] ^ 14);
  assign w647[8] = |(datain[279:276] ^ 1);
  assign w647[9] = |(datain[275:272] ^ 15);
  assign w647[10] = |(datain[271:268] ^ 11);
  assign w647[11] = |(datain[267:264] ^ 11);
  assign w647[12] = |(datain[263:260] ^ 4);
  assign w647[13] = |(datain[259:256] ^ 9);
  assign w647[14] = |(datain[255:252] ^ 1);
  assign w647[15] = |(datain[251:248] ^ 0);
  assign w647[16] = |(datain[247:244] ^ 4);
  assign w647[17] = |(datain[243:240] ^ 3);
  assign w647[18] = |(datain[239:236] ^ 3);
  assign w647[19] = |(datain[235:232] ^ 1);
  assign w647[20] = |(datain[231:228] ^ 5);
  assign w647[21] = |(datain[227:224] ^ 7);
  assign w647[22] = |(datain[223:220] ^ 6);
  assign w647[23] = |(datain[219:216] ^ 13);
  assign w647[24] = |(datain[215:212] ^ 3);
  assign w647[25] = |(datain[211:208] ^ 1);
  assign w647[26] = |(datain[207:204] ^ 4);
  assign w647[27] = |(datain[203:200] ^ 15);
  assign w647[28] = |(datain[199:196] ^ 6);
  assign w647[29] = |(datain[195:192] ^ 13);
  assign w647[30] = |(datain[191:188] ^ 3);
  assign w647[31] = |(datain[187:184] ^ 1);
  assign w647[32] = |(datain[183:180] ^ 5);
  assign w647[33] = |(datain[179:176] ^ 15);
  assign w647[34] = |(datain[175:172] ^ 6);
  assign w647[35] = |(datain[171:168] ^ 13);
  assign w647[36] = |(datain[167:164] ^ 14);
  assign w647[37] = |(datain[163:160] ^ 2);
  assign w647[38] = |(datain[159:156] ^ 15);
  assign w647[39] = |(datain[155:152] ^ 4);
  assign comp[647] = ~(|w647);
  wire [48-1:0] w648;
  assign w648[0] = |(datain[311:308] ^ 4);
  assign w648[1] = |(datain[307:304] ^ 0);
  assign w648[2] = |(datain[303:300] ^ 11);
  assign w648[3] = |(datain[299:296] ^ 9);
  assign w648[4] = |(datain[295:292] ^ 13);
  assign w648[5] = |(datain[291:288] ^ 1);
  assign w648[6] = |(datain[287:284] ^ 0);
  assign w648[7] = |(datain[283:280] ^ 0);
  assign w648[8] = |(datain[279:276] ^ 9);
  assign w648[9] = |(datain[275:272] ^ 9);
  assign w648[10] = |(datain[271:268] ^ 12);
  assign w648[11] = |(datain[267:264] ^ 13);
  assign w648[12] = |(datain[263:260] ^ 2);
  assign w648[13] = |(datain[259:256] ^ 1);
  assign w648[14] = |(datain[255:252] ^ 11);
  assign w648[15] = |(datain[251:248] ^ 8);
  assign w648[16] = |(datain[247:244] ^ 0);
  assign w648[17] = |(datain[243:240] ^ 0);
  assign w648[18] = |(datain[239:236] ^ 4);
  assign w648[19] = |(datain[235:232] ^ 2);
  assign w648[20] = |(datain[231:228] ^ 3);
  assign w648[21] = |(datain[227:224] ^ 3);
  assign w648[22] = |(datain[223:220] ^ 12);
  assign w648[23] = |(datain[219:216] ^ 9);
  assign w648[24] = |(datain[215:212] ^ 12);
  assign w648[25] = |(datain[211:208] ^ 13);
  assign w648[26] = |(datain[207:204] ^ 2);
  assign w648[27] = |(datain[203:200] ^ 1);
  assign w648[28] = |(datain[199:196] ^ 11);
  assign w648[29] = |(datain[195:192] ^ 4);
  assign w648[30] = |(datain[191:188] ^ 4);
  assign w648[31] = |(datain[187:184] ^ 0);
  assign w648[32] = |(datain[183:180] ^ 11);
  assign w648[33] = |(datain[179:176] ^ 1);
  assign w648[34] = |(datain[175:172] ^ 1);
  assign w648[35] = |(datain[171:168] ^ 8);
  assign w648[36] = |(datain[167:164] ^ 11);
  assign w648[37] = |(datain[163:160] ^ 10);
  assign w648[38] = |(datain[159:156] ^ 13);
  assign w648[39] = |(datain[155:152] ^ 1);
  assign w648[40] = |(datain[151:148] ^ 0);
  assign w648[41] = |(datain[147:144] ^ 0);
  assign w648[42] = |(datain[143:140] ^ 12);
  assign w648[43] = |(datain[139:136] ^ 13);
  assign w648[44] = |(datain[135:132] ^ 2);
  assign w648[45] = |(datain[131:128] ^ 1);
  assign w648[46] = |(datain[127:124] ^ 11);
  assign w648[47] = |(datain[123:120] ^ 4);
  assign comp[648] = ~(|w648);
  wire [76-1:0] w649;
  assign w649[0] = |(datain[311:308] ^ 12);
  assign w649[1] = |(datain[307:304] ^ 0);
  assign w649[2] = |(datain[303:300] ^ 0);
  assign w649[3] = |(datain[299:296] ^ 1);
  assign w649[4] = |(datain[295:292] ^ 11);
  assign w649[5] = |(datain[291:288] ^ 8);
  assign w649[6] = |(datain[287:284] ^ 11);
  assign w649[7] = |(datain[283:280] ^ 4);
  assign w649[8] = |(datain[279:276] ^ 4);
  assign w649[9] = |(datain[275:272] ^ 0);
  assign w649[10] = |(datain[271:268] ^ 11);
  assign w649[11] = |(datain[267:264] ^ 9);
  assign w649[12] = |(datain[263:260] ^ 14);
  assign w649[13] = |(datain[259:256] ^ 7);
  assign w649[14] = |(datain[255:252] ^ 0);
  assign w649[15] = |(datain[251:248] ^ 0);
  assign w649[16] = |(datain[247:244] ^ 11);
  assign w649[17] = |(datain[243:240] ^ 10);
  assign w649[18] = |(datain[239:236] ^ 0);
  assign w649[19] = |(datain[235:232] ^ 0);
  assign w649[20] = |(datain[231:228] ^ 0);
  assign w649[21] = |(datain[227:224] ^ 1);
  assign w649[22] = |(datain[223:220] ^ 12);
  assign w649[23] = |(datain[219:216] ^ 13);
  assign w649[24] = |(datain[215:212] ^ 2);
  assign w649[25] = |(datain[211:208] ^ 1);
  assign w649[26] = |(datain[207:204] ^ 11);
  assign w649[27] = |(datain[203:200] ^ 8);
  assign w649[28] = |(datain[199:196] ^ 0);
  assign w649[29] = |(datain[195:192] ^ 0);
  assign w649[30] = |(datain[191:188] ^ 4);
  assign w649[31] = |(datain[187:184] ^ 2);
  assign w649[32] = |(datain[183:180] ^ 3);
  assign w649[33] = |(datain[179:176] ^ 3);
  assign w649[34] = |(datain[175:172] ^ 12);
  assign w649[35] = |(datain[171:168] ^ 9);
  assign w649[36] = |(datain[167:164] ^ 3);
  assign w649[37] = |(datain[163:160] ^ 3);
  assign w649[38] = |(datain[159:156] ^ 13);
  assign w649[39] = |(datain[155:152] ^ 2);
  assign w649[40] = |(datain[151:148] ^ 12);
  assign w649[41] = |(datain[147:144] ^ 13);
  assign w649[42] = |(datain[143:140] ^ 2);
  assign w649[43] = |(datain[139:136] ^ 1);
  assign w649[44] = |(datain[135:132] ^ 11);
  assign w649[45] = |(datain[131:128] ^ 4);
  assign w649[46] = |(datain[127:124] ^ 4);
  assign w649[47] = |(datain[123:120] ^ 0);
  assign w649[48] = |(datain[119:116] ^ 11);
  assign w649[49] = |(datain[115:112] ^ 9);
  assign w649[50] = |(datain[111:108] ^ 0);
  assign w649[51] = |(datain[107:104] ^ 4);
  assign w649[52] = |(datain[103:100] ^ 0);
  assign w649[53] = |(datain[99:96] ^ 0);
  assign w649[54] = |(datain[95:92] ^ 11);
  assign w649[55] = |(datain[91:88] ^ 10);
  assign w649[56] = |(datain[87:84] ^ 0);
  assign w649[57] = |(datain[83:80] ^ 0);
  assign w649[58] = |(datain[79:76] ^ 0);
  assign w649[59] = |(datain[75:72] ^ 1);
  assign w649[60] = |(datain[71:68] ^ 12);
  assign w649[61] = |(datain[67:64] ^ 13);
  assign w649[62] = |(datain[63:60] ^ 2);
  assign w649[63] = |(datain[59:56] ^ 1);
  assign w649[64] = |(datain[55:52] ^ 5);
  assign w649[65] = |(datain[51:48] ^ 10);
  assign w649[66] = |(datain[47:44] ^ 5);
  assign w649[67] = |(datain[43:40] ^ 9);
  assign w649[68] = |(datain[39:36] ^ 5);
  assign w649[69] = |(datain[35:32] ^ 8);
  assign w649[70] = |(datain[31:28] ^ 4);
  assign w649[71] = |(datain[27:24] ^ 0);
  assign w649[72] = |(datain[23:20] ^ 12);
  assign w649[73] = |(datain[19:16] ^ 13);
  assign w649[74] = |(datain[15:12] ^ 2);
  assign w649[75] = |(datain[11:8] ^ 1);
  assign comp[649] = ~(|w649);
  wire [32-1:0] w650;
  assign w650[0] = |(datain[311:308] ^ 8);
  assign w650[1] = |(datain[307:304] ^ 12);
  assign w650[2] = |(datain[303:300] ^ 0);
  assign w650[3] = |(datain[299:296] ^ 6);
  assign w650[4] = |(datain[295:292] ^ 5);
  assign w650[5] = |(datain[291:288] ^ 11);
  assign w650[6] = |(datain[287:284] ^ 0);
  assign w650[7] = |(datain[283:280] ^ 1);
  assign w650[8] = |(datain[279:276] ^ 8);
  assign w650[9] = |(datain[275:272] ^ 12);
  assign w650[10] = |(datain[271:268] ^ 12);
  assign w650[11] = |(datain[267:264] ^ 8);
  assign w650[12] = |(datain[263:260] ^ 8);
  assign w650[13] = |(datain[259:256] ^ 14);
  assign w650[14] = |(datain[255:252] ^ 13);
  assign w650[15] = |(datain[251:248] ^ 8);
  assign w650[16] = |(datain[247:244] ^ 11);
  assign w650[17] = |(datain[243:240] ^ 8);
  assign w650[18] = |(datain[239:236] ^ 2);
  assign w650[19] = |(datain[235:232] ^ 1);
  assign w650[20] = |(datain[231:228] ^ 2);
  assign w650[21] = |(datain[227:224] ^ 5);
  assign w650[22] = |(datain[223:220] ^ 11);
  assign w650[23] = |(datain[219:216] ^ 10);
  assign w650[24] = |(datain[215:212] ^ 9);
  assign w650[25] = |(datain[211:208] ^ 4);
  assign w650[26] = |(datain[207:204] ^ 0);
  assign w650[27] = |(datain[203:200] ^ 1);
  assign w650[28] = |(datain[199:196] ^ 12);
  assign w650[29] = |(datain[195:192] ^ 13);
  assign w650[30] = |(datain[191:188] ^ 2);
  assign w650[31] = |(datain[187:184] ^ 1);
  assign comp[650] = ~(|w650);
  wire [74-1:0] w651;
  assign w651[0] = |(datain[311:308] ^ 5);
  assign w651[1] = |(datain[307:304] ^ 11);
  assign w651[2] = |(datain[303:300] ^ 8);
  assign w651[3] = |(datain[299:296] ^ 1);
  assign w651[4] = |(datain[295:292] ^ 14);
  assign w651[5] = |(datain[291:288] ^ 11);
  assign w651[6] = |(datain[287:284] ^ 0);
  assign w651[7] = |(datain[283:280] ^ 6);
  assign w651[8] = |(datain[279:276] ^ 0);
  assign w651[9] = |(datain[275:272] ^ 1);
  assign w651[10] = |(datain[271:268] ^ 14);
  assign w651[11] = |(datain[267:264] ^ 4);
  assign w651[12] = |(datain[263:260] ^ 2);
  assign w651[13] = |(datain[259:256] ^ 1);
  assign w651[14] = |(datain[255:252] ^ 10);
  assign w651[15] = |(datain[251:248] ^ 2);
  assign w651[16] = |(datain[247:244] ^ 15);
  assign w651[17] = |(datain[243:240] ^ 15);
  assign w651[18] = |(datain[239:236] ^ 0);
  assign w651[19] = |(datain[235:232] ^ 0);
  assign w651[20] = |(datain[231:228] ^ 11);
  assign w651[21] = |(datain[227:224] ^ 0);
  assign w651[22] = |(datain[223:220] ^ 15);
  assign w651[23] = |(datain[219:216] ^ 14);
  assign w651[24] = |(datain[215:212] ^ 14);
  assign w651[25] = |(datain[211:208] ^ 6);
  assign w651[26] = |(datain[207:204] ^ 2);
  assign w651[27] = |(datain[203:200] ^ 1);
  assign w651[28] = |(datain[199:196] ^ 11);
  assign w651[29] = |(datain[195:192] ^ 14);
  assign w651[30] = |(datain[191:188] ^ 0);
  assign w651[31] = |(datain[187:184] ^ 1);
  assign w651[32] = |(datain[183:180] ^ 0);
  assign w651[33] = |(datain[179:176] ^ 1);
  assign w651[34] = |(datain[175:172] ^ 8);
  assign w651[35] = |(datain[171:168] ^ 9);
  assign w651[36] = |(datain[167:164] ^ 15);
  assign w651[37] = |(datain[163:160] ^ 7);
  assign w651[38] = |(datain[159:156] ^ 15);
  assign w651[39] = |(datain[155:152] ^ 11);
  assign w651[40] = |(datain[151:148] ^ 15);
  assign w651[41] = |(datain[147:144] ^ 4);
  assign w651[42] = |(datain[143:140] ^ 3);
  assign w651[43] = |(datain[139:136] ^ 3);
  assign w651[44] = |(datain[135:132] ^ 12);
  assign w651[45] = |(datain[131:128] ^ 0);
  assign w651[46] = |(datain[127:124] ^ 8);
  assign w651[47] = |(datain[123:120] ^ 14);
  assign w651[48] = |(datain[119:116] ^ 13);
  assign w651[49] = |(datain[115:112] ^ 0);
  assign w651[50] = |(datain[111:108] ^ 8);
  assign w651[51] = |(datain[107:104] ^ 9);
  assign w651[52] = |(datain[103:100] ^ 12);
  assign w651[53] = |(datain[99:96] ^ 4);
  assign w651[54] = |(datain[95:92] ^ 8);
  assign w651[55] = |(datain[91:88] ^ 12);
  assign w651[56] = |(datain[87:84] ^ 12);
  assign w651[57] = |(datain[83:80] ^ 8);
  assign w651[58] = |(datain[79:76] ^ 8);
  assign w651[59] = |(datain[75:72] ^ 14);
  assign w651[60] = |(datain[71:68] ^ 13);
  assign w651[61] = |(datain[67:64] ^ 8);
  assign w651[62] = |(datain[63:60] ^ 8);
  assign w651[63] = |(datain[59:56] ^ 15);
  assign w651[64] = |(datain[55:52] ^ 0);
  assign w651[65] = |(datain[51:48] ^ 4);
  assign w651[66] = |(datain[47:44] ^ 15);
  assign w651[67] = |(datain[43:40] ^ 15);
  assign w651[68] = |(datain[39:36] ^ 3);
  assign w651[69] = |(datain[35:32] ^ 5);
  assign w651[70] = |(datain[31:28] ^ 5);
  assign w651[71] = |(datain[27:24] ^ 8);
  assign w651[72] = |(datain[23:20] ^ 8);
  assign w651[73] = |(datain[19:16] ^ 3);
  assign comp[651] = ~(|w651);
  wire [60-1:0] w652;
  assign w652[0] = |(datain[311:308] ^ 0);
  assign w652[1] = |(datain[307:304] ^ 4);
  assign w652[2] = |(datain[303:300] ^ 11);
  assign w652[3] = |(datain[299:296] ^ 10);
  assign w652[4] = |(datain[295:292] ^ 0);
  assign w652[5] = |(datain[291:288] ^ 0);
  assign w652[6] = |(datain[287:284] ^ 0);
  assign w652[7] = |(datain[283:280] ^ 1);
  assign w652[8] = |(datain[279:276] ^ 11);
  assign w652[9] = |(datain[275:272] ^ 4);
  assign w652[10] = |(datain[271:268] ^ 4);
  assign w652[11] = |(datain[267:264] ^ 0);
  assign w652[12] = |(datain[263:260] ^ 12);
  assign w652[13] = |(datain[259:256] ^ 13);
  assign w652[14] = |(datain[255:252] ^ 2);
  assign w652[15] = |(datain[251:248] ^ 1);
  assign w652[16] = |(datain[247:244] ^ 11);
  assign w652[17] = |(datain[243:240] ^ 8);
  assign w652[18] = |(datain[239:236] ^ 0);
  assign w652[19] = |(datain[235:232] ^ 0);
  assign w652[20] = |(datain[231:228] ^ 4);
  assign w652[21] = |(datain[227:224] ^ 2);
  assign w652[22] = |(datain[223:220] ^ 3);
  assign w652[23] = |(datain[219:216] ^ 3);
  assign w652[24] = |(datain[215:212] ^ 12);
  assign w652[25] = |(datain[211:208] ^ 9);
  assign w652[26] = |(datain[207:204] ^ 3);
  assign w652[27] = |(datain[203:200] ^ 3);
  assign w652[28] = |(datain[199:196] ^ 13);
  assign w652[29] = |(datain[195:192] ^ 2);
  assign w652[30] = |(datain[191:188] ^ 12);
  assign w652[31] = |(datain[187:184] ^ 13);
  assign w652[32] = |(datain[183:180] ^ 2);
  assign w652[33] = |(datain[179:176] ^ 1);
  assign w652[34] = |(datain[175:172] ^ 11);
  assign w652[35] = |(datain[171:168] ^ 4);
  assign w652[36] = |(datain[167:164] ^ 4);
  assign w652[37] = |(datain[163:160] ^ 0);
  assign w652[38] = |(datain[159:156] ^ 11);
  assign w652[39] = |(datain[155:152] ^ 9);
  assign w652[40] = |(datain[151:148] ^ 0);
  assign w652[41] = |(datain[147:144] ^ 7);
  assign w652[42] = |(datain[143:140] ^ 0);
  assign w652[43] = |(datain[139:136] ^ 0);
  assign w652[44] = |(datain[135:132] ^ 11);
  assign w652[45] = |(datain[131:128] ^ 10);
  assign w652[46] = |(datain[127:124] ^ 0);
  assign w652[47] = |(datain[123:120] ^ 0);
  assign w652[48] = |(datain[119:116] ^ 0);
  assign w652[49] = |(datain[115:112] ^ 1);
  assign w652[50] = |(datain[111:108] ^ 12);
  assign w652[51] = |(datain[107:104] ^ 13);
  assign w652[52] = |(datain[103:100] ^ 2);
  assign w652[53] = |(datain[99:96] ^ 1);
  assign w652[54] = |(datain[95:92] ^ 11);
  assign w652[55] = |(datain[91:88] ^ 8);
  assign w652[56] = |(datain[87:84] ^ 0);
  assign w652[57] = |(datain[83:80] ^ 2);
  assign w652[58] = |(datain[79:76] ^ 4);
  assign w652[59] = |(datain[75:72] ^ 2);
  assign comp[652] = ~(|w652);
  wire [44-1:0] w653;
  assign w653[0] = |(datain[311:308] ^ 3);
  assign w653[1] = |(datain[307:304] ^ 3);
  assign w653[2] = |(datain[303:300] ^ 12);
  assign w653[3] = |(datain[299:296] ^ 9);
  assign w653[4] = |(datain[295:292] ^ 12);
  assign w653[5] = |(datain[291:288] ^ 13);
  assign w653[6] = |(datain[287:284] ^ 2);
  assign w653[7] = |(datain[283:280] ^ 1);
  assign w653[8] = |(datain[279:276] ^ 8);
  assign w653[9] = |(datain[275:272] ^ 11);
  assign w653[10] = |(datain[271:268] ^ 13);
  assign w653[11] = |(datain[267:264] ^ 8);
  assign w653[12] = |(datain[263:260] ^ 11);
  assign w653[13] = |(datain[259:256] ^ 4);
  assign w653[14] = |(datain[255:252] ^ 4);
  assign w653[15] = |(datain[251:248] ^ 0);
  assign w653[16] = |(datain[247:244] ^ 11);
  assign w653[17] = |(datain[243:240] ^ 9);
  assign w653[18] = |(datain[239:236] ^ 11);
  assign w653[19] = |(datain[235:232] ^ 12);
  assign w653[20] = |(datain[231:228] ^ 0);
  assign w653[21] = |(datain[227:224] ^ 2);
  assign w653[22] = |(datain[223:220] ^ 8);
  assign w653[23] = |(datain[219:216] ^ 13);
  assign w653[24] = |(datain[215:212] ^ 9);
  assign w653[25] = |(datain[211:208] ^ 6);
  assign w653[26] = |(datain[207:204] ^ 8);
  assign w653[27] = |(datain[203:200] ^ 11);
  assign w653[28] = |(datain[199:196] ^ 0);
  assign w653[29] = |(datain[195:192] ^ 1);
  assign w653[30] = |(datain[191:188] ^ 12);
  assign w653[31] = |(datain[187:184] ^ 13);
  assign w653[32] = |(datain[183:180] ^ 2);
  assign w653[33] = |(datain[179:176] ^ 1);
  assign w653[34] = |(datain[175:172] ^ 11);
  assign w653[35] = |(datain[171:168] ^ 4);
  assign w653[36] = |(datain[167:164] ^ 3);
  assign w653[37] = |(datain[163:160] ^ 14);
  assign w653[38] = |(datain[159:156] ^ 12);
  assign w653[39] = |(datain[155:152] ^ 13);
  assign w653[40] = |(datain[151:148] ^ 2);
  assign w653[41] = |(datain[147:144] ^ 1);
  assign w653[42] = |(datain[143:140] ^ 12);
  assign w653[43] = |(datain[139:136] ^ 3);
  assign comp[653] = ~(|w653);
  wire [42-1:0] w654;
  assign w654[0] = |(datain[311:308] ^ 9);
  assign w654[1] = |(datain[307:304] ^ 11);
  assign w654[2] = |(datain[303:300] ^ 0);
  assign w654[3] = |(datain[299:296] ^ 4);
  assign w654[4] = |(datain[295:292] ^ 11);
  assign w654[5] = |(datain[291:288] ^ 10);
  assign w654[6] = |(datain[287:284] ^ 0);
  assign w654[7] = |(datain[283:280] ^ 0);
  assign w654[8] = |(datain[279:276] ^ 0);
  assign w654[9] = |(datain[275:272] ^ 1);
  assign w654[10] = |(datain[271:268] ^ 12);
  assign w654[11] = |(datain[267:264] ^ 13);
  assign w654[12] = |(datain[263:260] ^ 2);
  assign w654[13] = |(datain[259:256] ^ 1);
  assign w654[14] = |(datain[255:252] ^ 11);
  assign w654[15] = |(datain[251:248] ^ 8);
  assign w654[16] = |(datain[247:244] ^ 0);
  assign w654[17] = |(datain[243:240] ^ 0);
  assign w654[18] = |(datain[239:236] ^ 4);
  assign w654[19] = |(datain[235:232] ^ 2);
  assign w654[20] = |(datain[231:228] ^ 3);
  assign w654[21] = |(datain[227:224] ^ 3);
  assign w654[22] = |(datain[223:220] ^ 12);
  assign w654[23] = |(datain[219:216] ^ 9);
  assign w654[24] = |(datain[215:212] ^ 3);
  assign w654[25] = |(datain[211:208] ^ 3);
  assign w654[26] = |(datain[207:204] ^ 13);
  assign w654[27] = |(datain[203:200] ^ 2);
  assign w654[28] = |(datain[199:196] ^ 12);
  assign w654[29] = |(datain[195:192] ^ 13);
  assign w654[30] = |(datain[191:188] ^ 2);
  assign w654[31] = |(datain[187:184] ^ 1);
  assign w654[32] = |(datain[183:180] ^ 12);
  assign w654[33] = |(datain[179:176] ^ 6);
  assign w654[34] = |(datain[175:172] ^ 0);
  assign w654[35] = |(datain[171:168] ^ 6);
  assign w654[36] = |(datain[167:164] ^ 4);
  assign w654[37] = |(datain[163:160] ^ 10);
  assign w654[38] = |(datain[159:156] ^ 0);
  assign w654[39] = |(datain[155:152] ^ 2);
  assign w654[40] = |(datain[151:148] ^ 5);
  assign w654[41] = |(datain[147:144] ^ 10);
  assign comp[654] = ~(|w654);
  wire [58-1:0] w655;
  assign w655[0] = |(datain[311:308] ^ 11);
  assign w655[1] = |(datain[307:304] ^ 4);
  assign w655[2] = |(datain[303:300] ^ 4);
  assign w655[3] = |(datain[299:296] ^ 0);
  assign w655[4] = |(datain[295:292] ^ 11);
  assign w655[5] = |(datain[291:288] ^ 1);
  assign w655[6] = |(datain[287:284] ^ 9);
  assign w655[7] = |(datain[283:280] ^ 8);
  assign w655[8] = |(datain[279:276] ^ 11);
  assign w655[9] = |(datain[275:272] ^ 6);
  assign w655[10] = |(datain[271:268] ^ 0);
  assign w655[11] = |(datain[267:264] ^ 1);
  assign w655[12] = |(datain[263:260] ^ 12);
  assign w655[13] = |(datain[259:256] ^ 13);
  assign w655[14] = |(datain[255:252] ^ 2);
  assign w655[15] = |(datain[251:248] ^ 1);
  assign w655[16] = |(datain[247:244] ^ 11);
  assign w655[17] = |(datain[243:240] ^ 8);
  assign w655[18] = |(datain[239:236] ^ 0);
  assign w655[19] = |(datain[235:232] ^ 0);
  assign w655[20] = |(datain[231:228] ^ 4);
  assign w655[21] = |(datain[227:224] ^ 2);
  assign w655[22] = |(datain[223:220] ^ 3);
  assign w655[23] = |(datain[219:216] ^ 3);
  assign w655[24] = |(datain[215:212] ^ 13);
  assign w655[25] = |(datain[211:208] ^ 2);
  assign w655[26] = |(datain[207:204] ^ 3);
  assign w655[27] = |(datain[203:200] ^ 3);
  assign w655[28] = |(datain[199:196] ^ 12);
  assign w655[29] = |(datain[195:192] ^ 9);
  assign w655[30] = |(datain[191:188] ^ 12);
  assign w655[31] = |(datain[187:184] ^ 13);
  assign w655[32] = |(datain[183:180] ^ 2);
  assign w655[33] = |(datain[179:176] ^ 1);
  assign w655[34] = |(datain[175:172] ^ 11);
  assign w655[35] = |(datain[171:168] ^ 4);
  assign w655[36] = |(datain[167:164] ^ 4);
  assign w655[37] = |(datain[163:160] ^ 0);
  assign w655[38] = |(datain[159:156] ^ 11);
  assign w655[39] = |(datain[155:152] ^ 6);
  assign w655[40] = |(datain[151:148] ^ 0);
  assign w655[41] = |(datain[147:144] ^ 1);
  assign w655[42] = |(datain[143:140] ^ 11);
  assign w655[43] = |(datain[139:136] ^ 1);
  assign w655[44] = |(datain[135:132] ^ 0);
  assign w655[45] = |(datain[131:128] ^ 4);
  assign w655[46] = |(datain[127:124] ^ 12);
  assign w655[47] = |(datain[123:120] ^ 13);
  assign w655[48] = |(datain[119:116] ^ 2);
  assign w655[49] = |(datain[115:112] ^ 1);
  assign w655[50] = |(datain[111:108] ^ 11);
  assign w655[51] = |(datain[107:104] ^ 4);
  assign w655[52] = |(datain[103:100] ^ 3);
  assign w655[53] = |(datain[99:96] ^ 14);
  assign w655[54] = |(datain[95:92] ^ 12);
  assign w655[55] = |(datain[91:88] ^ 13);
  assign w655[56] = |(datain[87:84] ^ 2);
  assign w655[57] = |(datain[83:80] ^ 1);
  assign comp[655] = ~(|w655);
  wire [60-1:0] w656;
  assign w656[0] = |(datain[311:308] ^ 0);
  assign w656[1] = |(datain[307:304] ^ 1);
  assign w656[2] = |(datain[303:300] ^ 11);
  assign w656[3] = |(datain[299:296] ^ 4);
  assign w656[4] = |(datain[295:292] ^ 4);
  assign w656[5] = |(datain[291:288] ^ 0);
  assign w656[6] = |(datain[287:284] ^ 11);
  assign w656[7] = |(datain[283:280] ^ 1);
  assign w656[8] = |(datain[279:276] ^ 9);
  assign w656[9] = |(datain[275:272] ^ 9);
  assign w656[10] = |(datain[271:268] ^ 11);
  assign w656[11] = |(datain[267:264] ^ 6);
  assign w656[12] = |(datain[263:260] ^ 0);
  assign w656[13] = |(datain[259:256] ^ 1);
  assign w656[14] = |(datain[255:252] ^ 12);
  assign w656[15] = |(datain[251:248] ^ 13);
  assign w656[16] = |(datain[247:244] ^ 2);
  assign w656[17] = |(datain[243:240] ^ 1);
  assign w656[18] = |(datain[239:236] ^ 11);
  assign w656[19] = |(datain[235:232] ^ 8);
  assign w656[20] = |(datain[231:228] ^ 0);
  assign w656[21] = |(datain[227:224] ^ 0);
  assign w656[22] = |(datain[223:220] ^ 4);
  assign w656[23] = |(datain[219:216] ^ 2);
  assign w656[24] = |(datain[215:212] ^ 3);
  assign w656[25] = |(datain[211:208] ^ 3);
  assign w656[26] = |(datain[207:204] ^ 13);
  assign w656[27] = |(datain[203:200] ^ 2);
  assign w656[28] = |(datain[199:196] ^ 3);
  assign w656[29] = |(datain[195:192] ^ 3);
  assign w656[30] = |(datain[191:188] ^ 12);
  assign w656[31] = |(datain[187:184] ^ 9);
  assign w656[32] = |(datain[183:180] ^ 12);
  assign w656[33] = |(datain[179:176] ^ 13);
  assign w656[34] = |(datain[175:172] ^ 2);
  assign w656[35] = |(datain[171:168] ^ 1);
  assign w656[36] = |(datain[167:164] ^ 11);
  assign w656[37] = |(datain[163:160] ^ 4);
  assign w656[38] = |(datain[159:156] ^ 4);
  assign w656[39] = |(datain[155:152] ^ 0);
  assign w656[40] = |(datain[151:148] ^ 11);
  assign w656[41] = |(datain[147:144] ^ 6);
  assign w656[42] = |(datain[143:140] ^ 0);
  assign w656[43] = |(datain[139:136] ^ 1);
  assign w656[44] = |(datain[135:132] ^ 11);
  assign w656[45] = |(datain[131:128] ^ 1);
  assign w656[46] = |(datain[127:124] ^ 0);
  assign w656[47] = |(datain[123:120] ^ 4);
  assign w656[48] = |(datain[119:116] ^ 12);
  assign w656[49] = |(datain[115:112] ^ 13);
  assign w656[50] = |(datain[111:108] ^ 2);
  assign w656[51] = |(datain[107:104] ^ 1);
  assign w656[52] = |(datain[103:100] ^ 11);
  assign w656[53] = |(datain[99:96] ^ 4);
  assign w656[54] = |(datain[95:92] ^ 3);
  assign w656[55] = |(datain[91:88] ^ 14);
  assign w656[56] = |(datain[87:84] ^ 12);
  assign w656[57] = |(datain[83:80] ^ 13);
  assign w656[58] = |(datain[79:76] ^ 2);
  assign w656[59] = |(datain[75:72] ^ 1);
  assign comp[656] = ~(|w656);
  wire [58-1:0] w657;
  assign w657[0] = |(datain[311:308] ^ 11);
  assign w657[1] = |(datain[307:304] ^ 4);
  assign w657[2] = |(datain[303:300] ^ 4);
  assign w657[3] = |(datain[299:296] ^ 0);
  assign w657[4] = |(datain[295:292] ^ 11);
  assign w657[5] = |(datain[291:288] ^ 1);
  assign w657[6] = |(datain[287:284] ^ 9);
  assign w657[7] = |(datain[283:280] ^ 11);
  assign w657[8] = |(datain[279:276] ^ 11);
  assign w657[9] = |(datain[275:272] ^ 6);
  assign w657[10] = |(datain[271:268] ^ 0);
  assign w657[11] = |(datain[267:264] ^ 1);
  assign w657[12] = |(datain[263:260] ^ 12);
  assign w657[13] = |(datain[259:256] ^ 13);
  assign w657[14] = |(datain[255:252] ^ 2);
  assign w657[15] = |(datain[251:248] ^ 1);
  assign w657[16] = |(datain[247:244] ^ 11);
  assign w657[17] = |(datain[243:240] ^ 8);
  assign w657[18] = |(datain[239:236] ^ 0);
  assign w657[19] = |(datain[235:232] ^ 0);
  assign w657[20] = |(datain[231:228] ^ 4);
  assign w657[21] = |(datain[227:224] ^ 2);
  assign w657[22] = |(datain[223:220] ^ 3);
  assign w657[23] = |(datain[219:216] ^ 3);
  assign w657[24] = |(datain[215:212] ^ 13);
  assign w657[25] = |(datain[211:208] ^ 2);
  assign w657[26] = |(datain[207:204] ^ 3);
  assign w657[27] = |(datain[203:200] ^ 3);
  assign w657[28] = |(datain[199:196] ^ 12);
  assign w657[29] = |(datain[195:192] ^ 9);
  assign w657[30] = |(datain[191:188] ^ 12);
  assign w657[31] = |(datain[187:184] ^ 13);
  assign w657[32] = |(datain[183:180] ^ 2);
  assign w657[33] = |(datain[179:176] ^ 1);
  assign w657[34] = |(datain[175:172] ^ 11);
  assign w657[35] = |(datain[171:168] ^ 4);
  assign w657[36] = |(datain[167:164] ^ 4);
  assign w657[37] = |(datain[163:160] ^ 0);
  assign w657[38] = |(datain[159:156] ^ 11);
  assign w657[39] = |(datain[155:152] ^ 6);
  assign w657[40] = |(datain[151:148] ^ 0);
  assign w657[41] = |(datain[147:144] ^ 1);
  assign w657[42] = |(datain[143:140] ^ 11);
  assign w657[43] = |(datain[139:136] ^ 1);
  assign w657[44] = |(datain[135:132] ^ 0);
  assign w657[45] = |(datain[131:128] ^ 4);
  assign w657[46] = |(datain[127:124] ^ 12);
  assign w657[47] = |(datain[123:120] ^ 13);
  assign w657[48] = |(datain[119:116] ^ 2);
  assign w657[49] = |(datain[115:112] ^ 1);
  assign w657[50] = |(datain[111:108] ^ 11);
  assign w657[51] = |(datain[107:104] ^ 4);
  assign w657[52] = |(datain[103:100] ^ 3);
  assign w657[53] = |(datain[99:96] ^ 14);
  assign w657[54] = |(datain[95:92] ^ 12);
  assign w657[55] = |(datain[91:88] ^ 13);
  assign w657[56] = |(datain[87:84] ^ 2);
  assign w657[57] = |(datain[83:80] ^ 1);
  assign comp[657] = ~(|w657);
  wire [46-1:0] w658;
  assign w658[0] = |(datain[311:308] ^ 0);
  assign w658[1] = |(datain[307:304] ^ 2);
  assign w658[2] = |(datain[303:300] ^ 3);
  assign w658[3] = |(datain[299:296] ^ 13);
  assign w658[4] = |(datain[295:292] ^ 11);
  assign w658[5] = |(datain[291:288] ^ 10);
  assign w658[6] = |(datain[287:284] ^ 9);
  assign w658[7] = |(datain[283:280] ^ 14);
  assign w658[8] = |(datain[279:276] ^ 0);
  assign w658[9] = |(datain[275:272] ^ 0);
  assign w658[10] = |(datain[271:268] ^ 12);
  assign w658[11] = |(datain[267:264] ^ 13);
  assign w658[12] = |(datain[263:260] ^ 2);
  assign w658[13] = |(datain[259:256] ^ 1);
  assign w658[14] = |(datain[255:252] ^ 8);
  assign w658[15] = |(datain[251:248] ^ 11);
  assign w658[16] = |(datain[247:244] ^ 13);
  assign w658[17] = |(datain[243:240] ^ 8);
  assign w658[18] = |(datain[239:236] ^ 11);
  assign w658[19] = |(datain[235:232] ^ 9);
  assign w658[20] = |(datain[231:228] ^ 0);
  assign w658[21] = |(datain[227:224] ^ 5);
  assign w658[22] = |(datain[223:220] ^ 0);
  assign w658[23] = |(datain[219:216] ^ 0);
  assign w658[24] = |(datain[215:212] ^ 8);
  assign w658[25] = |(datain[211:208] ^ 13);
  assign w658[26] = |(datain[207:204] ^ 9);
  assign w658[27] = |(datain[203:200] ^ 6);
  assign w658[28] = |(datain[199:196] ^ 2);
  assign w658[29] = |(datain[195:192] ^ 1);
  assign w658[30] = |(datain[191:188] ^ 0);
  assign w658[31] = |(datain[187:184] ^ 1);
  assign w658[32] = |(datain[183:180] ^ 11);
  assign w658[33] = |(datain[179:176] ^ 4);
  assign w658[34] = |(datain[175:172] ^ 3);
  assign w658[35] = |(datain[171:168] ^ 15);
  assign w658[36] = |(datain[167:164] ^ 12);
  assign w658[37] = |(datain[163:160] ^ 13);
  assign w658[38] = |(datain[159:156] ^ 2);
  assign w658[39] = |(datain[155:152] ^ 1);
  assign w658[40] = |(datain[151:148] ^ 8);
  assign w658[41] = |(datain[147:144] ^ 9);
  assign w658[42] = |(datain[143:140] ^ 13);
  assign w658[43] = |(datain[139:136] ^ 6);
  assign w658[44] = |(datain[135:132] ^ 10);
  assign w658[45] = |(datain[131:128] ^ 13);
  assign comp[658] = ~(|w658);
  wire [60-1:0] w659;
  assign w659[0] = |(datain[311:308] ^ 10);
  assign w659[1] = |(datain[307:304] ^ 3);
  assign w659[2] = |(datain[303:300] ^ 0);
  assign w659[3] = |(datain[299:296] ^ 5);
  assign w659[4] = |(datain[295:292] ^ 0);
  assign w659[5] = |(datain[291:288] ^ 1);
  assign w659[6] = |(datain[287:284] ^ 11);
  assign w659[7] = |(datain[283:280] ^ 4);
  assign w659[8] = |(datain[279:276] ^ 4);
  assign w659[9] = |(datain[275:272] ^ 0);
  assign w659[10] = |(datain[271:268] ^ 11);
  assign w659[11] = |(datain[267:264] ^ 9);
  assign w659[12] = |(datain[263:260] ^ 11);
  assign w659[13] = |(datain[259:256] ^ 11);
  assign w659[14] = |(datain[255:252] ^ 0);
  assign w659[15] = |(datain[251:248] ^ 0);
  assign w659[16] = |(datain[247:244] ^ 11);
  assign w659[17] = |(datain[243:240] ^ 10);
  assign w659[18] = |(datain[239:236] ^ 0);
  assign w659[19] = |(datain[235:232] ^ 0);
  assign w659[20] = |(datain[231:228] ^ 0);
  assign w659[21] = |(datain[227:224] ^ 1);
  assign w659[22] = |(datain[223:220] ^ 12);
  assign w659[23] = |(datain[219:216] ^ 13);
  assign w659[24] = |(datain[215:212] ^ 2);
  assign w659[25] = |(datain[211:208] ^ 1);
  assign w659[26] = |(datain[207:204] ^ 11);
  assign w659[27] = |(datain[203:200] ^ 8);
  assign w659[28] = |(datain[199:196] ^ 0);
  assign w659[29] = |(datain[195:192] ^ 0);
  assign w659[30] = |(datain[191:188] ^ 4);
  assign w659[31] = |(datain[187:184] ^ 2);
  assign w659[32] = |(datain[183:180] ^ 3);
  assign w659[33] = |(datain[179:176] ^ 3);
  assign w659[34] = |(datain[175:172] ^ 13);
  assign w659[35] = |(datain[171:168] ^ 2);
  assign w659[36] = |(datain[167:164] ^ 3);
  assign w659[37] = |(datain[163:160] ^ 3);
  assign w659[38] = |(datain[159:156] ^ 12);
  assign w659[39] = |(datain[155:152] ^ 9);
  assign w659[40] = |(datain[151:148] ^ 12);
  assign w659[41] = |(datain[147:144] ^ 13);
  assign w659[42] = |(datain[143:140] ^ 2);
  assign w659[43] = |(datain[139:136] ^ 1);
  assign w659[44] = |(datain[135:132] ^ 11);
  assign w659[45] = |(datain[131:128] ^ 4);
  assign w659[46] = |(datain[127:124] ^ 4);
  assign w659[47] = |(datain[123:120] ^ 0);
  assign w659[48] = |(datain[119:116] ^ 11);
  assign w659[49] = |(datain[115:112] ^ 6);
  assign w659[50] = |(datain[111:108] ^ 0);
  assign w659[51] = |(datain[107:104] ^ 1);
  assign w659[52] = |(datain[103:100] ^ 11);
  assign w659[53] = |(datain[99:96] ^ 1);
  assign w659[54] = |(datain[95:92] ^ 0);
  assign w659[55] = |(datain[91:88] ^ 4);
  assign w659[56] = |(datain[87:84] ^ 12);
  assign w659[57] = |(datain[83:80] ^ 13);
  assign w659[58] = |(datain[79:76] ^ 2);
  assign w659[59] = |(datain[75:72] ^ 1);
  assign comp[659] = ~(|w659);
  wire [42-1:0] w660;
  assign w660[0] = |(datain[311:308] ^ 13);
  assign w660[1] = |(datain[307:304] ^ 5);
  assign w660[2] = |(datain[303:300] ^ 12);
  assign w660[3] = |(datain[299:296] ^ 13);
  assign w660[4] = |(datain[295:292] ^ 2);
  assign w660[5] = |(datain[291:288] ^ 1);
  assign w660[6] = |(datain[287:284] ^ 11);
  assign w660[7] = |(datain[283:280] ^ 8);
  assign w660[8] = |(datain[279:276] ^ 0);
  assign w660[9] = |(datain[275:272] ^ 0);
  assign w660[10] = |(datain[271:268] ^ 4);
  assign w660[11] = |(datain[267:264] ^ 2);
  assign w660[12] = |(datain[263:260] ^ 2);
  assign w660[13] = |(datain[259:256] ^ 11);
  assign w660[14] = |(datain[255:252] ^ 12);
  assign w660[15] = |(datain[251:248] ^ 9);
  assign w660[16] = |(datain[247:244] ^ 2);
  assign w660[17] = |(datain[243:240] ^ 11);
  assign w660[18] = |(datain[239:236] ^ 13);
  assign w660[19] = |(datain[235:232] ^ 2);
  assign w660[20] = |(datain[231:228] ^ 12);
  assign w660[21] = |(datain[227:224] ^ 13);
  assign w660[22] = |(datain[223:220] ^ 2);
  assign w660[23] = |(datain[219:216] ^ 1);
  assign w660[24] = |(datain[215:212] ^ 11);
  assign w660[25] = |(datain[211:208] ^ 4);
  assign w660[26] = |(datain[207:204] ^ 4);
  assign w660[27] = |(datain[203:200] ^ 0);
  assign w660[28] = |(datain[199:196] ^ 11);
  assign w660[29] = |(datain[195:192] ^ 1);
  assign w660[30] = |(datain[191:188] ^ 0);
  assign w660[31] = |(datain[187:184] ^ 3);
  assign w660[32] = |(datain[183:180] ^ 11);
  assign w660[33] = |(datain[179:176] ^ 6);
  assign w660[34] = |(datain[175:172] ^ 0);
  assign w660[35] = |(datain[171:168] ^ 1);
  assign w660[36] = |(datain[167:164] ^ 12);
  assign w660[37] = |(datain[163:160] ^ 13);
  assign w660[38] = |(datain[159:156] ^ 2);
  assign w660[39] = |(datain[155:152] ^ 1);
  assign w660[40] = |(datain[151:148] ^ 5);
  assign w660[41] = |(datain[147:144] ^ 10);
  assign comp[660] = ~(|w660);
  wire [64-1:0] w661;
  assign w661[0] = |(datain[311:308] ^ 0);
  assign w661[1] = |(datain[307:304] ^ 2);
  assign w661[2] = |(datain[303:300] ^ 0);
  assign w661[3] = |(datain[299:296] ^ 1);
  assign w661[4] = |(datain[295:292] ^ 10);
  assign w661[5] = |(datain[291:288] ^ 3);
  assign w661[6] = |(datain[287:284] ^ 0);
  assign w661[7] = |(datain[283:280] ^ 5);
  assign w661[8] = |(datain[279:276] ^ 0);
  assign w661[9] = |(datain[275:272] ^ 1);
  assign w661[10] = |(datain[271:268] ^ 11);
  assign w661[11] = |(datain[267:264] ^ 4);
  assign w661[12] = |(datain[263:260] ^ 4);
  assign w661[13] = |(datain[259:256] ^ 0);
  assign w661[14] = |(datain[255:252] ^ 11);
  assign w661[15] = |(datain[251:248] ^ 9);
  assign w661[16] = |(datain[247:244] ^ 13);
  assign w661[17] = |(datain[243:240] ^ 7);
  assign w661[18] = |(datain[239:236] ^ 0);
  assign w661[19] = |(datain[235:232] ^ 0);
  assign w661[20] = |(datain[231:228] ^ 11);
  assign w661[21] = |(datain[227:224] ^ 10);
  assign w661[22] = |(datain[223:220] ^ 0);
  assign w661[23] = |(datain[219:216] ^ 0);
  assign w661[24] = |(datain[215:212] ^ 0);
  assign w661[25] = |(datain[211:208] ^ 1);
  assign w661[26] = |(datain[207:204] ^ 12);
  assign w661[27] = |(datain[203:200] ^ 13);
  assign w661[28] = |(datain[199:196] ^ 2);
  assign w661[29] = |(datain[195:192] ^ 1);
  assign w661[30] = |(datain[191:188] ^ 11);
  assign w661[31] = |(datain[187:184] ^ 8);
  assign w661[32] = |(datain[183:180] ^ 0);
  assign w661[33] = |(datain[179:176] ^ 0);
  assign w661[34] = |(datain[175:172] ^ 4);
  assign w661[35] = |(datain[171:168] ^ 2);
  assign w661[36] = |(datain[167:164] ^ 3);
  assign w661[37] = |(datain[163:160] ^ 3);
  assign w661[38] = |(datain[159:156] ^ 13);
  assign w661[39] = |(datain[155:152] ^ 2);
  assign w661[40] = |(datain[151:148] ^ 3);
  assign w661[41] = |(datain[147:144] ^ 3);
  assign w661[42] = |(datain[143:140] ^ 12);
  assign w661[43] = |(datain[139:136] ^ 9);
  assign w661[44] = |(datain[135:132] ^ 12);
  assign w661[45] = |(datain[131:128] ^ 13);
  assign w661[46] = |(datain[127:124] ^ 2);
  assign w661[47] = |(datain[123:120] ^ 1);
  assign w661[48] = |(datain[119:116] ^ 11);
  assign w661[49] = |(datain[115:112] ^ 4);
  assign w661[50] = |(datain[111:108] ^ 4);
  assign w661[51] = |(datain[107:104] ^ 0);
  assign w661[52] = |(datain[103:100] ^ 11);
  assign w661[53] = |(datain[99:96] ^ 6);
  assign w661[54] = |(datain[95:92] ^ 0);
  assign w661[55] = |(datain[91:88] ^ 1);
  assign w661[56] = |(datain[87:84] ^ 11);
  assign w661[57] = |(datain[83:80] ^ 1);
  assign w661[58] = |(datain[79:76] ^ 0);
  assign w661[59] = |(datain[75:72] ^ 4);
  assign w661[60] = |(datain[71:68] ^ 12);
  assign w661[61] = |(datain[67:64] ^ 13);
  assign w661[62] = |(datain[63:60] ^ 2);
  assign w661[63] = |(datain[59:56] ^ 1);
  assign comp[661] = ~(|w661);
  wire [46-1:0] w662;
  assign w662[0] = |(datain[311:308] ^ 4);
  assign w662[1] = |(datain[307:304] ^ 0);
  assign w662[2] = |(datain[303:300] ^ 11);
  assign w662[3] = |(datain[299:296] ^ 1);
  assign w662[4] = |(datain[295:292] ^ 13);
  assign w662[5] = |(datain[291:288] ^ 9);
  assign w662[6] = |(datain[287:284] ^ 12);
  assign w662[7] = |(datain[283:280] ^ 13);
  assign w662[8] = |(datain[279:276] ^ 2);
  assign w662[9] = |(datain[275:272] ^ 1);
  assign w662[10] = |(datain[271:268] ^ 11);
  assign w662[11] = |(datain[267:264] ^ 8);
  assign w662[12] = |(datain[263:260] ^ 0);
  assign w662[13] = |(datain[259:256] ^ 0);
  assign w662[14] = |(datain[255:252] ^ 4);
  assign w662[15] = |(datain[251:248] ^ 2);
  assign w662[16] = |(datain[247:244] ^ 2);
  assign w662[17] = |(datain[243:240] ^ 11);
  assign w662[18] = |(datain[239:236] ^ 12);
  assign w662[19] = |(datain[235:232] ^ 9);
  assign w662[20] = |(datain[231:228] ^ 2);
  assign w662[21] = |(datain[227:224] ^ 11);
  assign w662[22] = |(datain[223:220] ^ 13);
  assign w662[23] = |(datain[219:216] ^ 2);
  assign w662[24] = |(datain[215:212] ^ 12);
  assign w662[25] = |(datain[211:208] ^ 13);
  assign w662[26] = |(datain[207:204] ^ 2);
  assign w662[27] = |(datain[203:200] ^ 1);
  assign w662[28] = |(datain[199:196] ^ 11);
  assign w662[29] = |(datain[195:192] ^ 4);
  assign w662[30] = |(datain[191:188] ^ 4);
  assign w662[31] = |(datain[187:184] ^ 0);
  assign w662[32] = |(datain[183:180] ^ 11);
  assign w662[33] = |(datain[179:176] ^ 1);
  assign w662[34] = |(datain[175:172] ^ 0);
  assign w662[35] = |(datain[171:168] ^ 3);
  assign w662[36] = |(datain[167:164] ^ 11);
  assign w662[37] = |(datain[163:160] ^ 6);
  assign w662[38] = |(datain[159:156] ^ 0);
  assign w662[39] = |(datain[155:152] ^ 1);
  assign w662[40] = |(datain[151:148] ^ 12);
  assign w662[41] = |(datain[147:144] ^ 13);
  assign w662[42] = |(datain[143:140] ^ 2);
  assign w662[43] = |(datain[139:136] ^ 1);
  assign w662[44] = |(datain[135:132] ^ 5);
  assign w662[45] = |(datain[131:128] ^ 10);
  assign comp[662] = ~(|w662);
  wire [42-1:0] w663;
  assign w663[0] = |(datain[311:308] ^ 13);
  assign w663[1] = |(datain[307:304] ^ 13);
  assign w663[2] = |(datain[303:300] ^ 0);
  assign w663[3] = |(datain[299:296] ^ 0);
  assign w663[4] = |(datain[295:292] ^ 12);
  assign w663[5] = |(datain[291:288] ^ 13);
  assign w663[6] = |(datain[287:284] ^ 2);
  assign w663[7] = |(datain[283:280] ^ 1);
  assign w663[8] = |(datain[279:276] ^ 11);
  assign w663[9] = |(datain[275:272] ^ 8);
  assign w663[10] = |(datain[271:268] ^ 0);
  assign w663[11] = |(datain[267:264] ^ 0);
  assign w663[12] = |(datain[263:260] ^ 4);
  assign w663[13] = |(datain[259:256] ^ 2);
  assign w663[14] = |(datain[255:252] ^ 2);
  assign w663[15] = |(datain[251:248] ^ 11);
  assign w663[16] = |(datain[247:244] ^ 12);
  assign w663[17] = |(datain[243:240] ^ 9);
  assign w663[18] = |(datain[239:236] ^ 2);
  assign w663[19] = |(datain[235:232] ^ 11);
  assign w663[20] = |(datain[231:228] ^ 13);
  assign w663[21] = |(datain[227:224] ^ 2);
  assign w663[22] = |(datain[223:220] ^ 12);
  assign w663[23] = |(datain[219:216] ^ 13);
  assign w663[24] = |(datain[215:212] ^ 2);
  assign w663[25] = |(datain[211:208] ^ 1);
  assign w663[26] = |(datain[207:204] ^ 11);
  assign w663[27] = |(datain[203:200] ^ 4);
  assign w663[28] = |(datain[199:196] ^ 4);
  assign w663[29] = |(datain[195:192] ^ 0);
  assign w663[30] = |(datain[191:188] ^ 11);
  assign w663[31] = |(datain[187:184] ^ 1);
  assign w663[32] = |(datain[183:180] ^ 0);
  assign w663[33] = |(datain[179:176] ^ 3);
  assign w663[34] = |(datain[175:172] ^ 11);
  assign w663[35] = |(datain[171:168] ^ 6);
  assign w663[36] = |(datain[167:164] ^ 0);
  assign w663[37] = |(datain[163:160] ^ 1);
  assign w663[38] = |(datain[159:156] ^ 12);
  assign w663[39] = |(datain[155:152] ^ 13);
  assign w663[40] = |(datain[151:148] ^ 2);
  assign w663[41] = |(datain[147:144] ^ 1);
  assign comp[663] = ~(|w663);
  wire [44-1:0] w664;
  assign w664[0] = |(datain[311:308] ^ 11);
  assign w664[1] = |(datain[307:304] ^ 9);
  assign w664[2] = |(datain[303:300] ^ 14);
  assign w664[3] = |(datain[299:296] ^ 5);
  assign w664[4] = |(datain[295:292] ^ 0);
  assign w664[5] = |(datain[291:288] ^ 0);
  assign w664[6] = |(datain[287:284] ^ 12);
  assign w664[7] = |(datain[283:280] ^ 13);
  assign w664[8] = |(datain[279:276] ^ 2);
  assign w664[9] = |(datain[275:272] ^ 1);
  assign w664[10] = |(datain[271:268] ^ 11);
  assign w664[11] = |(datain[267:264] ^ 8);
  assign w664[12] = |(datain[263:260] ^ 0);
  assign w664[13] = |(datain[259:256] ^ 0);
  assign w664[14] = |(datain[255:252] ^ 4);
  assign w664[15] = |(datain[251:248] ^ 2);
  assign w664[16] = |(datain[247:244] ^ 2);
  assign w664[17] = |(datain[243:240] ^ 11);
  assign w664[18] = |(datain[239:236] ^ 12);
  assign w664[19] = |(datain[235:232] ^ 9);
  assign w664[20] = |(datain[231:228] ^ 2);
  assign w664[21] = |(datain[227:224] ^ 11);
  assign w664[22] = |(datain[223:220] ^ 13);
  assign w664[23] = |(datain[219:216] ^ 2);
  assign w664[24] = |(datain[215:212] ^ 12);
  assign w664[25] = |(datain[211:208] ^ 13);
  assign w664[26] = |(datain[207:204] ^ 2);
  assign w664[27] = |(datain[203:200] ^ 1);
  assign w664[28] = |(datain[199:196] ^ 11);
  assign w664[29] = |(datain[195:192] ^ 4);
  assign w664[30] = |(datain[191:188] ^ 4);
  assign w664[31] = |(datain[187:184] ^ 0);
  assign w664[32] = |(datain[183:180] ^ 11);
  assign w664[33] = |(datain[179:176] ^ 1);
  assign w664[34] = |(datain[175:172] ^ 0);
  assign w664[35] = |(datain[171:168] ^ 3);
  assign w664[36] = |(datain[167:164] ^ 11);
  assign w664[37] = |(datain[163:160] ^ 6);
  assign w664[38] = |(datain[159:156] ^ 0);
  assign w664[39] = |(datain[155:152] ^ 1);
  assign w664[40] = |(datain[151:148] ^ 12);
  assign w664[41] = |(datain[147:144] ^ 13);
  assign w664[42] = |(datain[143:140] ^ 2);
  assign w664[43] = |(datain[139:136] ^ 1);
  assign comp[664] = ~(|w664);
  wire [56-1:0] w665;
  assign w665[0] = |(datain[311:308] ^ 11);
  assign w665[1] = |(datain[307:304] ^ 4);
  assign w665[2] = |(datain[303:300] ^ 4);
  assign w665[3] = |(datain[299:296] ^ 0);
  assign w665[4] = |(datain[295:292] ^ 11);
  assign w665[5] = |(datain[291:288] ^ 9);
  assign w665[6] = |(datain[287:284] ^ 3);
  assign w665[7] = |(datain[283:280] ^ 2);
  assign w665[8] = |(datain[279:276] ^ 0);
  assign w665[9] = |(datain[275:272] ^ 1);
  assign w665[10] = |(datain[271:268] ^ 12);
  assign w665[11] = |(datain[267:264] ^ 13);
  assign w665[12] = |(datain[263:260] ^ 2);
  assign w665[13] = |(datain[259:256] ^ 1);
  assign w665[14] = |(datain[255:252] ^ 11);
  assign w665[15] = |(datain[251:248] ^ 8);
  assign w665[16] = |(datain[247:244] ^ 0);
  assign w665[17] = |(datain[243:240] ^ 0);
  assign w665[18] = |(datain[239:236] ^ 4);
  assign w665[19] = |(datain[235:232] ^ 2);
  assign w665[20] = |(datain[231:228] ^ 3);
  assign w665[21] = |(datain[227:224] ^ 3);
  assign w665[22] = |(datain[223:220] ^ 13);
  assign w665[23] = |(datain[219:216] ^ 2);
  assign w665[24] = |(datain[215:212] ^ 3);
  assign w665[25] = |(datain[211:208] ^ 3);
  assign w665[26] = |(datain[207:204] ^ 12);
  assign w665[27] = |(datain[203:200] ^ 9);
  assign w665[28] = |(datain[199:196] ^ 12);
  assign w665[29] = |(datain[195:192] ^ 13);
  assign w665[30] = |(datain[191:188] ^ 2);
  assign w665[31] = |(datain[187:184] ^ 1);
  assign w665[32] = |(datain[183:180] ^ 11);
  assign w665[33] = |(datain[179:176] ^ 4);
  assign w665[34] = |(datain[175:172] ^ 4);
  assign w665[35] = |(datain[171:168] ^ 0);
  assign w665[36] = |(datain[167:164] ^ 11);
  assign w665[37] = |(datain[163:160] ^ 9);
  assign w665[38] = |(datain[159:156] ^ 0);
  assign w665[39] = |(datain[155:152] ^ 4);
  assign w665[40] = |(datain[151:148] ^ 0);
  assign w665[41] = |(datain[147:144] ^ 0);
  assign w665[42] = |(datain[143:140] ^ 11);
  assign w665[43] = |(datain[139:136] ^ 10);
  assign w665[44] = |(datain[135:132] ^ 5);
  assign w665[45] = |(datain[131:128] ^ 14);
  assign w665[46] = |(datain[127:124] ^ 0);
  assign w665[47] = |(datain[123:120] ^ 1);
  assign w665[48] = |(datain[119:116] ^ 12);
  assign w665[49] = |(datain[115:112] ^ 13);
  assign w665[50] = |(datain[111:108] ^ 2);
  assign w665[51] = |(datain[107:104] ^ 1);
  assign w665[52] = |(datain[103:100] ^ 5);
  assign w665[53] = |(datain[99:96] ^ 10);
  assign w665[54] = |(datain[95:92] ^ 5);
  assign w665[55] = |(datain[91:88] ^ 9);
  assign comp[665] = ~(|w665);
  wire [66-1:0] w666;
  assign w666[0] = |(datain[311:308] ^ 0);
  assign w666[1] = |(datain[307:304] ^ 6);
  assign w666[2] = |(datain[303:300] ^ 14);
  assign w666[3] = |(datain[299:296] ^ 15);
  assign w666[4] = |(datain[295:292] ^ 0);
  assign w666[5] = |(datain[291:288] ^ 1);
  assign w666[6] = |(datain[287:284] ^ 11);
  assign w666[7] = |(datain[283:280] ^ 8);
  assign w666[8] = |(datain[279:276] ^ 11);
  assign w666[9] = |(datain[275:272] ^ 4);
  assign w666[10] = |(datain[271:268] ^ 4);
  assign w666[11] = |(datain[267:264] ^ 0);
  assign w666[12] = |(datain[263:260] ^ 11);
  assign w666[13] = |(datain[259:256] ^ 9);
  assign w666[14] = |(datain[255:252] ^ 5);
  assign w666[15] = |(datain[251:248] ^ 2);
  assign w666[16] = |(datain[247:244] ^ 0);
  assign w666[17] = |(datain[243:240] ^ 1);
  assign w666[18] = |(datain[239:236] ^ 11);
  assign w666[19] = |(datain[235:232] ^ 10);
  assign w666[20] = |(datain[231:228] ^ 0);
  assign w666[21] = |(datain[227:224] ^ 0);
  assign w666[22] = |(datain[223:220] ^ 0);
  assign w666[23] = |(datain[219:216] ^ 1);
  assign w666[24] = |(datain[215:212] ^ 12);
  assign w666[25] = |(datain[211:208] ^ 13);
  assign w666[26] = |(datain[207:204] ^ 2);
  assign w666[27] = |(datain[203:200] ^ 1);
  assign w666[28] = |(datain[199:196] ^ 11);
  assign w666[29] = |(datain[195:192] ^ 8);
  assign w666[30] = |(datain[191:188] ^ 0);
  assign w666[31] = |(datain[187:184] ^ 0);
  assign w666[32] = |(datain[183:180] ^ 4);
  assign w666[33] = |(datain[179:176] ^ 2);
  assign w666[34] = |(datain[175:172] ^ 3);
  assign w666[35] = |(datain[171:168] ^ 3);
  assign w666[36] = |(datain[167:164] ^ 12);
  assign w666[37] = |(datain[163:160] ^ 9);
  assign w666[38] = |(datain[159:156] ^ 3);
  assign w666[39] = |(datain[155:152] ^ 3);
  assign w666[40] = |(datain[151:148] ^ 13);
  assign w666[41] = |(datain[147:144] ^ 2);
  assign w666[42] = |(datain[143:140] ^ 12);
  assign w666[43] = |(datain[139:136] ^ 13);
  assign w666[44] = |(datain[135:132] ^ 2);
  assign w666[45] = |(datain[131:128] ^ 1);
  assign w666[46] = |(datain[127:124] ^ 11);
  assign w666[47] = |(datain[123:120] ^ 9);
  assign w666[48] = |(datain[119:116] ^ 0);
  assign w666[49] = |(datain[115:112] ^ 3);
  assign w666[50] = |(datain[111:108] ^ 0);
  assign w666[51] = |(datain[107:104] ^ 0);
  assign w666[52] = |(datain[103:100] ^ 11);
  assign w666[53] = |(datain[99:96] ^ 10);
  assign w666[54] = |(datain[95:92] ^ 0);
  assign w666[55] = |(datain[91:88] ^ 0);
  assign w666[56] = |(datain[87:84] ^ 0);
  assign w666[57] = |(datain[83:80] ^ 1);
  assign w666[58] = |(datain[79:76] ^ 11);
  assign w666[59] = |(datain[75:72] ^ 4);
  assign w666[60] = |(datain[71:68] ^ 4);
  assign w666[61] = |(datain[67:64] ^ 0);
  assign w666[62] = |(datain[63:60] ^ 12);
  assign w666[63] = |(datain[59:56] ^ 13);
  assign w666[64] = |(datain[55:52] ^ 2);
  assign w666[65] = |(datain[51:48] ^ 1);
  assign comp[666] = ~(|w666);
  wire [58-1:0] w667;
  assign w667[0] = |(datain[311:308] ^ 4);
  assign w667[1] = |(datain[307:304] ^ 0);
  assign w667[2] = |(datain[303:300] ^ 11);
  assign w667[3] = |(datain[299:296] ^ 10);
  assign w667[4] = |(datain[295:292] ^ 0);
  assign w667[5] = |(datain[291:288] ^ 0);
  assign w667[6] = |(datain[287:284] ^ 0);
  assign w667[7] = |(datain[283:280] ^ 1);
  assign w667[8] = |(datain[279:276] ^ 11);
  assign w667[9] = |(datain[275:272] ^ 9);
  assign w667[10] = |(datain[271:268] ^ 7);
  assign w667[11] = |(datain[267:264] ^ 1);
  assign w667[12] = |(datain[263:260] ^ 0);
  assign w667[13] = |(datain[259:256] ^ 1);
  assign w667[14] = |(datain[255:252] ^ 0);
  assign w667[15] = |(datain[251:248] ^ 3);
  assign w667[16] = |(datain[247:244] ^ 1);
  assign w667[17] = |(datain[243:240] ^ 6);
  assign w667[18] = |(datain[239:236] ^ 0);
  assign w667[19] = |(datain[235:232] ^ 1);
  assign w667[20] = |(datain[231:228] ^ 0);
  assign w667[21] = |(datain[227:224] ^ 1);
  assign w667[22] = |(datain[223:220] ^ 12);
  assign w667[23] = |(datain[219:216] ^ 13);
  assign w667[24] = |(datain[215:212] ^ 2);
  assign w667[25] = |(datain[211:208] ^ 1);
  assign w667[26] = |(datain[207:204] ^ 11);
  assign w667[27] = |(datain[203:200] ^ 9);
  assign w667[28] = |(datain[199:196] ^ 3);
  assign w667[29] = |(datain[195:192] ^ 12);
  assign w667[30] = |(datain[191:188] ^ 0);
  assign w667[31] = |(datain[187:184] ^ 0);
  assign w667[32] = |(datain[183:180] ^ 11);
  assign w667[33] = |(datain[179:176] ^ 14);
  assign w667[34] = |(datain[175:172] ^ 3);
  assign w667[35] = |(datain[171:168] ^ 4);
  assign w667[36] = |(datain[167:164] ^ 0);
  assign w667[37] = |(datain[163:160] ^ 2);
  assign w667[38] = |(datain[159:156] ^ 0);
  assign w667[39] = |(datain[155:152] ^ 3);
  assign w667[40] = |(datain[151:148] ^ 3);
  assign w667[41] = |(datain[147:144] ^ 6);
  assign w667[42] = |(datain[143:140] ^ 0);
  assign w667[43] = |(datain[139:136] ^ 1);
  assign w667[44] = |(datain[135:132] ^ 0);
  assign w667[45] = |(datain[131:128] ^ 1);
  assign w667[46] = |(datain[127:124] ^ 8);
  assign w667[47] = |(datain[123:120] ^ 0);
  assign w667[48] = |(datain[119:116] ^ 3);
  assign w667[49] = |(datain[115:112] ^ 4);
  assign w667[50] = |(datain[111:108] ^ 0);
  assign w667[51] = |(datain[107:104] ^ 1);
  assign w667[52] = |(datain[103:100] ^ 4);
  assign w667[53] = |(datain[99:96] ^ 6);
  assign w667[54] = |(datain[95:92] ^ 14);
  assign w667[55] = |(datain[91:88] ^ 2);
  assign w667[56] = |(datain[87:84] ^ 15);
  assign w667[57] = |(datain[83:80] ^ 10);
  assign comp[667] = ~(|w667);
  wire [56-1:0] w668;
  assign w668[0] = |(datain[311:308] ^ 4);
  assign w668[1] = |(datain[307:304] ^ 0);
  assign w668[2] = |(datain[303:300] ^ 11);
  assign w668[3] = |(datain[299:296] ^ 9);
  assign w668[4] = |(datain[295:292] ^ 7);
  assign w668[5] = |(datain[291:288] ^ 9);
  assign w668[6] = |(datain[287:284] ^ 0);
  assign w668[7] = |(datain[283:280] ^ 1);
  assign w668[8] = |(datain[279:276] ^ 11);
  assign w668[9] = |(datain[275:272] ^ 10);
  assign w668[10] = |(datain[271:268] ^ 0);
  assign w668[11] = |(datain[267:264] ^ 0);
  assign w668[12] = |(datain[263:260] ^ 0);
  assign w668[13] = |(datain[259:256] ^ 0);
  assign w668[14] = |(datain[255:252] ^ 12);
  assign w668[15] = |(datain[251:248] ^ 13);
  assign w668[16] = |(datain[247:244] ^ 2);
  assign w668[17] = |(datain[243:240] ^ 1);
  assign w668[18] = |(datain[239:236] ^ 11);
  assign w668[19] = |(datain[235:232] ^ 8);
  assign w668[20] = |(datain[231:228] ^ 0);
  assign w668[21] = |(datain[227:224] ^ 0);
  assign w668[22] = |(datain[223:220] ^ 4);
  assign w668[23] = |(datain[219:216] ^ 2);
  assign w668[24] = |(datain[215:212] ^ 3);
  assign w668[25] = |(datain[211:208] ^ 3);
  assign w668[26] = |(datain[207:204] ^ 12);
  assign w668[27] = |(datain[203:200] ^ 9);
  assign w668[28] = |(datain[199:196] ^ 3);
  assign w668[29] = |(datain[195:192] ^ 3);
  assign w668[30] = |(datain[191:188] ^ 13);
  assign w668[31] = |(datain[187:184] ^ 2);
  assign w668[32] = |(datain[183:180] ^ 12);
  assign w668[33] = |(datain[179:176] ^ 13);
  assign w668[34] = |(datain[175:172] ^ 2);
  assign w668[35] = |(datain[171:168] ^ 1);
  assign w668[36] = |(datain[167:164] ^ 11);
  assign w668[37] = |(datain[163:160] ^ 9);
  assign w668[38] = |(datain[159:156] ^ 0);
  assign w668[39] = |(datain[155:152] ^ 3);
  assign w668[40] = |(datain[151:148] ^ 0);
  assign w668[41] = |(datain[147:144] ^ 0);
  assign w668[42] = |(datain[143:140] ^ 11);
  assign w668[43] = |(datain[139:136] ^ 10);
  assign w668[44] = |(datain[135:132] ^ 0);
  assign w668[45] = |(datain[131:128] ^ 0);
  assign w668[46] = |(datain[127:124] ^ 0);
  assign w668[47] = |(datain[123:120] ^ 0);
  assign w668[48] = |(datain[119:116] ^ 11);
  assign w668[49] = |(datain[115:112] ^ 4);
  assign w668[50] = |(datain[111:108] ^ 4);
  assign w668[51] = |(datain[107:104] ^ 0);
  assign w668[52] = |(datain[103:100] ^ 12);
  assign w668[53] = |(datain[99:96] ^ 13);
  assign w668[54] = |(datain[95:92] ^ 2);
  assign w668[55] = |(datain[91:88] ^ 1);
  assign comp[668] = ~(|w668);
  wire [58-1:0] w669;
  assign w669[0] = |(datain[311:308] ^ 11);
  assign w669[1] = |(datain[307:304] ^ 9);
  assign w669[2] = |(datain[303:300] ^ 3);
  assign w669[3] = |(datain[299:296] ^ 8);
  assign w669[4] = |(datain[295:292] ^ 0);
  assign w669[5] = |(datain[291:288] ^ 15);
  assign w669[6] = |(datain[287:284] ^ 11);
  assign w669[7] = |(datain[283:280] ^ 10);
  assign w669[8] = |(datain[279:276] ^ 0);
  assign w669[9] = |(datain[275:272] ^ 0);
  assign w669[10] = |(datain[271:268] ^ 0);
  assign w669[11] = |(datain[267:264] ^ 1);
  assign w669[12] = |(datain[263:260] ^ 12);
  assign w669[13] = |(datain[259:256] ^ 13);
  assign w669[14] = |(datain[255:252] ^ 2);
  assign w669[15] = |(datain[251:248] ^ 1);
  assign w669[16] = |(datain[247:244] ^ 11);
  assign w669[17] = |(datain[243:240] ^ 8);
  assign w669[18] = |(datain[239:236] ^ 0);
  assign w669[19] = |(datain[235:232] ^ 0);
  assign w669[20] = |(datain[231:228] ^ 4);
  assign w669[21] = |(datain[227:224] ^ 2);
  assign w669[22] = |(datain[223:220] ^ 3);
  assign w669[23] = |(datain[219:216] ^ 3);
  assign w669[24] = |(datain[215:212] ^ 13);
  assign w669[25] = |(datain[211:208] ^ 2);
  assign w669[26] = |(datain[207:204] ^ 3);
  assign w669[27] = |(datain[203:200] ^ 3);
  assign w669[28] = |(datain[199:196] ^ 12);
  assign w669[29] = |(datain[195:192] ^ 9);
  assign w669[30] = |(datain[191:188] ^ 12);
  assign w669[31] = |(datain[187:184] ^ 13);
  assign w669[32] = |(datain[183:180] ^ 2);
  assign w669[33] = |(datain[179:176] ^ 1);
  assign w669[34] = |(datain[175:172] ^ 11);
  assign w669[35] = |(datain[171:168] ^ 4);
  assign w669[36] = |(datain[167:164] ^ 4);
  assign w669[37] = |(datain[163:160] ^ 0);
  assign w669[38] = |(datain[159:156] ^ 11);
  assign w669[39] = |(datain[155:152] ^ 9);
  assign w669[40] = |(datain[151:148] ^ 0);
  assign w669[41] = |(datain[147:144] ^ 4);
  assign w669[42] = |(datain[143:140] ^ 0);
  assign w669[43] = |(datain[139:136] ^ 0);
  assign w669[44] = |(datain[135:132] ^ 11);
  assign w669[45] = |(datain[131:128] ^ 10);
  assign w669[46] = |(datain[127:124] ^ 0);
  assign w669[47] = |(datain[123:120] ^ 0);
  assign w669[48] = |(datain[119:116] ^ 0);
  assign w669[49] = |(datain[115:112] ^ 1);
  assign w669[50] = |(datain[111:108] ^ 12);
  assign w669[51] = |(datain[107:104] ^ 13);
  assign w669[52] = |(datain[103:100] ^ 2);
  assign w669[53] = |(datain[99:96] ^ 1);
  assign w669[54] = |(datain[95:92] ^ 5);
  assign w669[55] = |(datain[91:88] ^ 9);
  assign w669[56] = |(datain[87:84] ^ 5);
  assign w669[57] = |(datain[83:80] ^ 10);
  assign comp[669] = ~(|w669);
  wire [58-1:0] w670;
  assign w670[0] = |(datain[311:308] ^ 0);
  assign w670[1] = |(datain[307:304] ^ 1);
  assign w670[2] = |(datain[303:300] ^ 11);
  assign w670[3] = |(datain[299:296] ^ 4);
  assign w670[4] = |(datain[295:292] ^ 4);
  assign w670[5] = |(datain[291:288] ^ 0);
  assign w670[6] = |(datain[287:284] ^ 11);
  assign w670[7] = |(datain[283:280] ^ 9);
  assign w670[8] = |(datain[279:276] ^ 14);
  assign w670[9] = |(datain[275:272] ^ 2);
  assign w670[10] = |(datain[271:268] ^ 0);
  assign w670[11] = |(datain[267:264] ^ 1);
  assign w670[12] = |(datain[263:260] ^ 12);
  assign w670[13] = |(datain[259:256] ^ 13);
  assign w670[14] = |(datain[255:252] ^ 2);
  assign w670[15] = |(datain[251:248] ^ 1);
  assign w670[16] = |(datain[247:244] ^ 11);
  assign w670[17] = |(datain[243:240] ^ 8);
  assign w670[18] = |(datain[239:236] ^ 0);
  assign w670[19] = |(datain[235:232] ^ 0);
  assign w670[20] = |(datain[231:228] ^ 4);
  assign w670[21] = |(datain[227:224] ^ 2);
  assign w670[22] = |(datain[223:220] ^ 2);
  assign w670[23] = |(datain[219:216] ^ 11);
  assign w670[24] = |(datain[215:212] ^ 13);
  assign w670[25] = |(datain[211:208] ^ 2);
  assign w670[26] = |(datain[207:204] ^ 2);
  assign w670[27] = |(datain[203:200] ^ 11);
  assign w670[28] = |(datain[199:196] ^ 12);
  assign w670[29] = |(datain[195:192] ^ 9);
  assign w670[30] = |(datain[191:188] ^ 12);
  assign w670[31] = |(datain[187:184] ^ 13);
  assign w670[32] = |(datain[183:180] ^ 2);
  assign w670[33] = |(datain[179:176] ^ 1);
  assign w670[34] = |(datain[175:172] ^ 11);
  assign w670[35] = |(datain[171:168] ^ 4);
  assign w670[36] = |(datain[167:164] ^ 4);
  assign w670[37] = |(datain[163:160] ^ 0);
  assign w670[38] = |(datain[159:156] ^ 11);
  assign w670[39] = |(datain[155:152] ^ 9);
  assign w670[40] = |(datain[151:148] ^ 0);
  assign w670[41] = |(datain[147:144] ^ 4);
  assign w670[42] = |(datain[143:140] ^ 0);
  assign w670[43] = |(datain[139:136] ^ 0);
  assign w670[44] = |(datain[135:132] ^ 11);
  assign w670[45] = |(datain[131:128] ^ 10);
  assign w670[46] = |(datain[127:124] ^ 7);
  assign w670[47] = |(datain[123:120] ^ 9);
  assign w670[48] = |(datain[119:116] ^ 0);
  assign w670[49] = |(datain[115:112] ^ 1);
  assign w670[50] = |(datain[111:108] ^ 12);
  assign w670[51] = |(datain[107:104] ^ 13);
  assign w670[52] = |(datain[103:100] ^ 2);
  assign w670[53] = |(datain[99:96] ^ 1);
  assign w670[54] = |(datain[95:92] ^ 5);
  assign w670[55] = |(datain[91:88] ^ 10);
  assign w670[56] = |(datain[87:84] ^ 5);
  assign w670[57] = |(datain[83:80] ^ 9);
  assign comp[670] = ~(|w670);
  wire [58-1:0] w671;
  assign w671[0] = |(datain[311:308] ^ 11);
  assign w671[1] = |(datain[307:304] ^ 10);
  assign w671[2] = |(datain[303:300] ^ 0);
  assign w671[3] = |(datain[299:296] ^ 0);
  assign w671[4] = |(datain[295:292] ^ 0);
  assign w671[5] = |(datain[291:288] ^ 1);
  assign w671[6] = |(datain[287:284] ^ 11);
  assign w671[7] = |(datain[283:280] ^ 4);
  assign w671[8] = |(datain[279:276] ^ 4);
  assign w671[9] = |(datain[275:272] ^ 0);
  assign w671[10] = |(datain[271:268] ^ 12);
  assign w671[11] = |(datain[267:264] ^ 13);
  assign w671[12] = |(datain[263:260] ^ 2);
  assign w671[13] = |(datain[259:256] ^ 1);
  assign w671[14] = |(datain[255:252] ^ 11);
  assign w671[15] = |(datain[251:248] ^ 8);
  assign w671[16] = |(datain[247:244] ^ 0);
  assign w671[17] = |(datain[243:240] ^ 0);
  assign w671[18] = |(datain[239:236] ^ 4);
  assign w671[19] = |(datain[235:232] ^ 2);
  assign w671[20] = |(datain[231:228] ^ 3);
  assign w671[21] = |(datain[227:224] ^ 3);
  assign w671[22] = |(datain[223:220] ^ 12);
  assign w671[23] = |(datain[219:216] ^ 9);
  assign w671[24] = |(datain[215:212] ^ 3);
  assign w671[25] = |(datain[211:208] ^ 3);
  assign w671[26] = |(datain[207:204] ^ 13);
  assign w671[27] = |(datain[203:200] ^ 2);
  assign w671[28] = |(datain[199:196] ^ 12);
  assign w671[29] = |(datain[195:192] ^ 13);
  assign w671[30] = |(datain[191:188] ^ 2);
  assign w671[31] = |(datain[187:184] ^ 1);
  assign w671[32] = |(datain[183:180] ^ 11);
  assign w671[33] = |(datain[179:176] ^ 4);
  assign w671[34] = |(datain[175:172] ^ 4);
  assign w671[35] = |(datain[171:168] ^ 0);
  assign w671[36] = |(datain[167:164] ^ 11);
  assign w671[37] = |(datain[163:160] ^ 9);
  assign w671[38] = |(datain[159:156] ^ 0);
  assign w671[39] = |(datain[155:152] ^ 7);
  assign w671[40] = |(datain[151:148] ^ 0);
  assign w671[41] = |(datain[147:144] ^ 0);
  assign w671[42] = |(datain[143:140] ^ 11);
  assign w671[43] = |(datain[139:136] ^ 10);
  assign w671[44] = |(datain[135:132] ^ 0);
  assign w671[45] = |(datain[131:128] ^ 0);
  assign w671[46] = |(datain[127:124] ^ 0);
  assign w671[47] = |(datain[123:120] ^ 1);
  assign w671[48] = |(datain[119:116] ^ 12);
  assign w671[49] = |(datain[115:112] ^ 13);
  assign w671[50] = |(datain[111:108] ^ 2);
  assign w671[51] = |(datain[107:104] ^ 1);
  assign w671[52] = |(datain[103:100] ^ 11);
  assign w671[53] = |(datain[99:96] ^ 8);
  assign w671[54] = |(datain[95:92] ^ 0);
  assign w671[55] = |(datain[91:88] ^ 2);
  assign w671[56] = |(datain[87:84] ^ 4);
  assign w671[57] = |(datain[83:80] ^ 2);
  assign comp[671] = ~(|w671);
  wire [42-1:0] w672;
  assign w672[0] = |(datain[311:308] ^ 3);
  assign w672[1] = |(datain[307:304] ^ 3);
  assign w672[2] = |(datain[303:300] ^ 12);
  assign w672[3] = |(datain[299:296] ^ 9);
  assign w672[4] = |(datain[295:292] ^ 11);
  assign w672[5] = |(datain[291:288] ^ 10);
  assign w672[6] = |(datain[287:284] ^ 4);
  assign w672[7] = |(datain[283:280] ^ 4);
  assign w672[8] = |(datain[279:276] ^ 0);
  assign w672[9] = |(datain[275:272] ^ 2);
  assign w672[10] = |(datain[271:268] ^ 12);
  assign w672[11] = |(datain[267:264] ^ 13);
  assign w672[12] = |(datain[263:260] ^ 2);
  assign w672[13] = |(datain[259:256] ^ 1);
  assign w672[14] = |(datain[255:252] ^ 7);
  assign w672[15] = |(datain[251:248] ^ 2);
  assign w672[16] = |(datain[247:244] ^ 5);
  assign w672[17] = |(datain[243:240] ^ 12);
  assign w672[18] = |(datain[239:236] ^ 8);
  assign w672[19] = |(datain[235:232] ^ 11);
  assign w672[20] = |(datain[231:228] ^ 13);
  assign w672[21] = |(datain[227:224] ^ 8);
  assign w672[22] = |(datain[223:220] ^ 11);
  assign w672[23] = |(datain[219:216] ^ 10);
  assign w672[24] = |(datain[215:212] ^ 4);
  assign w672[25] = |(datain[211:208] ^ 5);
  assign w672[26] = |(datain[207:204] ^ 0);
  assign w672[27] = |(datain[203:200] ^ 1);
  assign w672[28] = |(datain[199:196] ^ 11);
  assign w672[29] = |(datain[195:192] ^ 9);
  assign w672[30] = |(datain[191:188] ^ 0);
  assign w672[31] = |(datain[187:184] ^ 5);
  assign w672[32] = |(datain[183:180] ^ 0);
  assign w672[33] = |(datain[179:176] ^ 0);
  assign w672[34] = |(datain[175:172] ^ 11);
  assign w672[35] = |(datain[171:168] ^ 4);
  assign w672[36] = |(datain[167:164] ^ 3);
  assign w672[37] = |(datain[163:160] ^ 15);
  assign w672[38] = |(datain[159:156] ^ 12);
  assign w672[39] = |(datain[155:152] ^ 13);
  assign w672[40] = |(datain[151:148] ^ 2);
  assign w672[41] = |(datain[147:144] ^ 1);
  assign comp[672] = ~(|w672);
  wire [46-1:0] w673;
  assign w673[0] = |(datain[311:308] ^ 4);
  assign w673[1] = |(datain[307:304] ^ 0);
  assign w673[2] = |(datain[303:300] ^ 11);
  assign w673[3] = |(datain[299:296] ^ 10);
  assign w673[4] = |(datain[295:292] ^ 0);
  assign w673[5] = |(datain[291:288] ^ 0);
  assign w673[6] = |(datain[287:284] ^ 0);
  assign w673[7] = |(datain[283:280] ^ 1);
  assign w673[8] = |(datain[279:276] ^ 11);
  assign w673[9] = |(datain[275:272] ^ 9);
  assign w673[10] = |(datain[271:268] ^ 4);
  assign w673[11] = |(datain[267:264] ^ 12);
  assign w673[12] = |(datain[263:260] ^ 0);
  assign w673[13] = |(datain[259:256] ^ 2);
  assign w673[14] = |(datain[255:252] ^ 12);
  assign w673[15] = |(datain[251:248] ^ 13);
  assign w673[16] = |(datain[247:244] ^ 2);
  assign w673[17] = |(datain[243:240] ^ 1);
  assign w673[18] = |(datain[239:236] ^ 11);
  assign w673[19] = |(datain[235:232] ^ 8);
  assign w673[20] = |(datain[231:228] ^ 0);
  assign w673[21] = |(datain[227:224] ^ 0);
  assign w673[22] = |(datain[223:220] ^ 4);
  assign w673[23] = |(datain[219:216] ^ 2);
  assign w673[24] = |(datain[215:212] ^ 3);
  assign w673[25] = |(datain[211:208] ^ 3);
  assign w673[26] = |(datain[207:204] ^ 13);
  assign w673[27] = |(datain[203:200] ^ 2);
  assign w673[28] = |(datain[199:196] ^ 3);
  assign w673[29] = |(datain[195:192] ^ 3);
  assign w673[30] = |(datain[191:188] ^ 12);
  assign w673[31] = |(datain[187:184] ^ 9);
  assign w673[32] = |(datain[183:180] ^ 12);
  assign w673[33] = |(datain[179:176] ^ 13);
  assign w673[34] = |(datain[175:172] ^ 2);
  assign w673[35] = |(datain[171:168] ^ 1);
  assign w673[36] = |(datain[167:164] ^ 11);
  assign w673[37] = |(datain[163:160] ^ 4);
  assign w673[38] = |(datain[159:156] ^ 4);
  assign w673[39] = |(datain[155:152] ^ 0);
  assign w673[40] = |(datain[151:148] ^ 11);
  assign w673[41] = |(datain[147:144] ^ 9);
  assign w673[42] = |(datain[143:140] ^ 0);
  assign w673[43] = |(datain[139:136] ^ 4);
  assign w673[44] = |(datain[135:132] ^ 0);
  assign w673[45] = |(datain[131:128] ^ 0);
  assign comp[673] = ~(|w673);
  wire [46-1:0] w674;
  assign w674[0] = |(datain[311:308] ^ 4);
  assign w674[1] = |(datain[307:304] ^ 0);
  assign w674[2] = |(datain[303:300] ^ 11);
  assign w674[3] = |(datain[299:296] ^ 9);
  assign w674[4] = |(datain[295:292] ^ 4);
  assign w674[5] = |(datain[291:288] ^ 15);
  assign w674[6] = |(datain[287:284] ^ 0);
  assign w674[7] = |(datain[283:280] ^ 2);
  assign w674[8] = |(datain[279:276] ^ 11);
  assign w674[9] = |(datain[275:272] ^ 10);
  assign w674[10] = |(datain[271:268] ^ 0);
  assign w674[11] = |(datain[267:264] ^ 0);
  assign w674[12] = |(datain[263:260] ^ 0);
  assign w674[13] = |(datain[259:256] ^ 1);
  assign w674[14] = |(datain[255:252] ^ 12);
  assign w674[15] = |(datain[251:248] ^ 13);
  assign w674[16] = |(datain[247:244] ^ 2);
  assign w674[17] = |(datain[243:240] ^ 1);
  assign w674[18] = |(datain[239:236] ^ 11);
  assign w674[19] = |(datain[235:232] ^ 8);
  assign w674[20] = |(datain[231:228] ^ 0);
  assign w674[21] = |(datain[227:224] ^ 0);
  assign w674[22] = |(datain[223:220] ^ 4);
  assign w674[23] = |(datain[219:216] ^ 2);
  assign w674[24] = |(datain[215:212] ^ 3);
  assign w674[25] = |(datain[211:208] ^ 3);
  assign w674[26] = |(datain[207:204] ^ 12);
  assign w674[27] = |(datain[203:200] ^ 9);
  assign w674[28] = |(datain[199:196] ^ 3);
  assign w674[29] = |(datain[195:192] ^ 3);
  assign w674[30] = |(datain[191:188] ^ 13);
  assign w674[31] = |(datain[187:184] ^ 2);
  assign w674[32] = |(datain[183:180] ^ 12);
  assign w674[33] = |(datain[179:176] ^ 13);
  assign w674[34] = |(datain[175:172] ^ 2);
  assign w674[35] = |(datain[171:168] ^ 1);
  assign w674[36] = |(datain[167:164] ^ 0);
  assign w674[37] = |(datain[163:160] ^ 14);
  assign w674[38] = |(datain[159:156] ^ 0);
  assign w674[39] = |(datain[155:152] ^ 14);
  assign w674[40] = |(datain[151:148] ^ 1);
  assign w674[41] = |(datain[147:144] ^ 15);
  assign w674[42] = |(datain[143:140] ^ 0);
  assign w674[43] = |(datain[139:136] ^ 7);
  assign w674[44] = |(datain[135:132] ^ 11);
  assign w674[45] = |(datain[131:128] ^ 10);
  assign comp[674] = ~(|w674);
  wire [42-1:0] w675;
  assign w675[0] = |(datain[311:308] ^ 12);
  assign w675[1] = |(datain[307:304] ^ 13);
  assign w675[2] = |(datain[303:300] ^ 2);
  assign w675[3] = |(datain[299:296] ^ 1);
  assign w675[4] = |(datain[295:292] ^ 7);
  assign w675[5] = |(datain[291:288] ^ 2);
  assign w675[6] = |(datain[287:284] ^ 6);
  assign w675[7] = |(datain[283:280] ^ 1);
  assign w675[8] = |(datain[279:276] ^ 8);
  assign w675[9] = |(datain[275:272] ^ 11);
  assign w675[10] = |(datain[271:268] ^ 13);
  assign w675[11] = |(datain[267:264] ^ 8);
  assign w675[12] = |(datain[263:260] ^ 0);
  assign w675[13] = |(datain[259:256] ^ 14);
  assign w675[14] = |(datain[255:252] ^ 0);
  assign w675[15] = |(datain[251:248] ^ 14);
  assign w675[16] = |(datain[247:244] ^ 0);
  assign w675[17] = |(datain[243:240] ^ 7);
  assign w675[18] = |(datain[239:236] ^ 1);
  assign w675[19] = |(datain[235:232] ^ 15);
  assign w675[20] = |(datain[231:228] ^ 11);
  assign w675[21] = |(datain[227:224] ^ 4);
  assign w675[22] = |(datain[223:220] ^ 3);
  assign w675[23] = |(datain[219:216] ^ 15);
  assign w675[24] = |(datain[215:212] ^ 11);
  assign w675[25] = |(datain[211:208] ^ 9);
  assign w675[26] = |(datain[207:204] ^ 0);
  assign w675[27] = |(datain[203:200] ^ 4);
  assign w675[28] = |(datain[199:196] ^ 0);
  assign w675[29] = |(datain[195:192] ^ 0);
  assign w675[30] = |(datain[191:188] ^ 11);
  assign w675[31] = |(datain[187:184] ^ 10);
  assign w675[32] = |(datain[183:180] ^ 7);
  assign w675[33] = |(datain[179:176] ^ 2);
  assign w675[34] = |(datain[175:172] ^ 0);
  assign w675[35] = |(datain[171:168] ^ 1);
  assign w675[36] = |(datain[167:164] ^ 12);
  assign w675[37] = |(datain[163:160] ^ 13);
  assign w675[38] = |(datain[159:156] ^ 2);
  assign w675[39] = |(datain[155:152] ^ 1);
  assign w675[40] = |(datain[151:148] ^ 8);
  assign w675[41] = |(datain[147:144] ^ 9);
  assign comp[675] = ~(|w675);
  wire [46-1:0] w676;
  assign w676[0] = |(datain[311:308] ^ 4);
  assign w676[1] = |(datain[307:304] ^ 0);
  assign w676[2] = |(datain[303:300] ^ 11);
  assign w676[3] = |(datain[299:296] ^ 9);
  assign w676[4] = |(datain[295:292] ^ 7);
  assign w676[5] = |(datain[291:288] ^ 11);
  assign w676[6] = |(datain[287:284] ^ 0);
  assign w676[7] = |(datain[283:280] ^ 2);
  assign w676[8] = |(datain[279:276] ^ 11);
  assign w676[9] = |(datain[275:272] ^ 10);
  assign w676[10] = |(datain[271:268] ^ 0);
  assign w676[11] = |(datain[267:264] ^ 0);
  assign w676[12] = |(datain[263:260] ^ 0);
  assign w676[13] = |(datain[259:256] ^ 1);
  assign w676[14] = |(datain[255:252] ^ 12);
  assign w676[15] = |(datain[251:248] ^ 13);
  assign w676[16] = |(datain[247:244] ^ 2);
  assign w676[17] = |(datain[243:240] ^ 1);
  assign w676[18] = |(datain[239:236] ^ 11);
  assign w676[19] = |(datain[235:232] ^ 8);
  assign w676[20] = |(datain[231:228] ^ 0);
  assign w676[21] = |(datain[227:224] ^ 0);
  assign w676[22] = |(datain[223:220] ^ 4);
  assign w676[23] = |(datain[219:216] ^ 2);
  assign w676[24] = |(datain[215:212] ^ 3);
  assign w676[25] = |(datain[211:208] ^ 3);
  assign w676[26] = |(datain[207:204] ^ 12);
  assign w676[27] = |(datain[203:200] ^ 9);
  assign w676[28] = |(datain[199:196] ^ 3);
  assign w676[29] = |(datain[195:192] ^ 3);
  assign w676[30] = |(datain[191:188] ^ 13);
  assign w676[31] = |(datain[187:184] ^ 2);
  assign w676[32] = |(datain[183:180] ^ 12);
  assign w676[33] = |(datain[179:176] ^ 13);
  assign w676[34] = |(datain[175:172] ^ 2);
  assign w676[35] = |(datain[171:168] ^ 1);
  assign w676[36] = |(datain[167:164] ^ 11);
  assign w676[37] = |(datain[163:160] ^ 4);
  assign w676[38] = |(datain[159:156] ^ 4);
  assign w676[39] = |(datain[155:152] ^ 0);
  assign w676[40] = |(datain[151:148] ^ 11);
  assign w676[41] = |(datain[147:144] ^ 9);
  assign w676[42] = |(datain[143:140] ^ 0);
  assign w676[43] = |(datain[139:136] ^ 4);
  assign w676[44] = |(datain[135:132] ^ 0);
  assign w676[45] = |(datain[131:128] ^ 0);
  assign comp[676] = ~(|w676);
  wire [44-1:0] w677;
  assign w677[0] = |(datain[311:308] ^ 11);
  assign w677[1] = |(datain[307:304] ^ 9);
  assign w677[2] = |(datain[303:300] ^ 13);
  assign w677[3] = |(datain[299:296] ^ 6);
  assign w677[4] = |(datain[295:292] ^ 0);
  assign w677[5] = |(datain[291:288] ^ 2);
  assign w677[6] = |(datain[287:284] ^ 12);
  assign w677[7] = |(datain[283:280] ^ 13);
  assign w677[8] = |(datain[279:276] ^ 2);
  assign w677[9] = |(datain[275:272] ^ 1);
  assign w677[10] = |(datain[271:268] ^ 11);
  assign w677[11] = |(datain[267:264] ^ 8);
  assign w677[12] = |(datain[263:260] ^ 0);
  assign w677[13] = |(datain[259:256] ^ 0);
  assign w677[14] = |(datain[255:252] ^ 4);
  assign w677[15] = |(datain[251:248] ^ 2);
  assign w677[16] = |(datain[247:244] ^ 3);
  assign w677[17] = |(datain[243:240] ^ 3);
  assign w677[18] = |(datain[239:236] ^ 13);
  assign w677[19] = |(datain[235:232] ^ 2);
  assign w677[20] = |(datain[231:228] ^ 3);
  assign w677[21] = |(datain[227:224] ^ 3);
  assign w677[22] = |(datain[223:220] ^ 12);
  assign w677[23] = |(datain[219:216] ^ 9);
  assign w677[24] = |(datain[215:212] ^ 12);
  assign w677[25] = |(datain[211:208] ^ 13);
  assign w677[26] = |(datain[207:204] ^ 2);
  assign w677[27] = |(datain[203:200] ^ 1);
  assign w677[28] = |(datain[199:196] ^ 11);
  assign w677[29] = |(datain[195:192] ^ 4);
  assign w677[30] = |(datain[191:188] ^ 4);
  assign w677[31] = |(datain[187:184] ^ 0);
  assign w677[32] = |(datain[183:180] ^ 11);
  assign w677[33] = |(datain[179:176] ^ 9);
  assign w677[34] = |(datain[175:172] ^ 0);
  assign w677[35] = |(datain[171:168] ^ 3);
  assign w677[36] = |(datain[167:164] ^ 0);
  assign w677[37] = |(datain[163:160] ^ 0);
  assign w677[38] = |(datain[159:156] ^ 11);
  assign w677[39] = |(datain[155:152] ^ 10);
  assign w677[40] = |(datain[151:148] ^ 0);
  assign w677[41] = |(datain[147:144] ^ 0);
  assign w677[42] = |(datain[143:140] ^ 0);
  assign w677[43] = |(datain[139:136] ^ 1);
  assign comp[677] = ~(|w677);
  wire [56-1:0] w678;
  assign w678[0] = |(datain[311:308] ^ 15);
  assign w678[1] = |(datain[307:304] ^ 10);
  assign w678[2] = |(datain[303:300] ^ 0);
  assign w678[3] = |(datain[299:296] ^ 2);
  assign w678[4] = |(datain[295:292] ^ 11);
  assign w678[5] = |(datain[291:288] ^ 10);
  assign w678[6] = |(datain[287:284] ^ 0);
  assign w678[7] = |(datain[283:280] ^ 0);
  assign w678[8] = |(datain[279:276] ^ 0);
  assign w678[9] = |(datain[275:272] ^ 1);
  assign w678[10] = |(datain[271:268] ^ 12);
  assign w678[11] = |(datain[267:264] ^ 13);
  assign w678[12] = |(datain[263:260] ^ 2);
  assign w678[13] = |(datain[259:256] ^ 1);
  assign w678[14] = |(datain[255:252] ^ 11);
  assign w678[15] = |(datain[251:248] ^ 8);
  assign w678[16] = |(datain[247:244] ^ 0);
  assign w678[17] = |(datain[243:240] ^ 0);
  assign w678[18] = |(datain[239:236] ^ 4);
  assign w678[19] = |(datain[235:232] ^ 2);
  assign w678[20] = |(datain[231:228] ^ 3);
  assign w678[21] = |(datain[227:224] ^ 3);
  assign w678[22] = |(datain[223:220] ^ 13);
  assign w678[23] = |(datain[219:216] ^ 2);
  assign w678[24] = |(datain[215:212] ^ 3);
  assign w678[25] = |(datain[211:208] ^ 3);
  assign w678[26] = |(datain[207:204] ^ 12);
  assign w678[27] = |(datain[203:200] ^ 9);
  assign w678[28] = |(datain[199:196] ^ 12);
  assign w678[29] = |(datain[195:192] ^ 13);
  assign w678[30] = |(datain[191:188] ^ 2);
  assign w678[31] = |(datain[187:184] ^ 1);
  assign w678[32] = |(datain[183:180] ^ 11);
  assign w678[33] = |(datain[179:176] ^ 4);
  assign w678[34] = |(datain[175:172] ^ 4);
  assign w678[35] = |(datain[171:168] ^ 0);
  assign w678[36] = |(datain[167:164] ^ 11);
  assign w678[37] = |(datain[163:160] ^ 9);
  assign w678[38] = |(datain[159:156] ^ 0);
  assign w678[39] = |(datain[155:152] ^ 4);
  assign w678[40] = |(datain[151:148] ^ 0);
  assign w678[41] = |(datain[147:144] ^ 0);
  assign w678[42] = |(datain[143:140] ^ 11);
  assign w678[43] = |(datain[139:136] ^ 10);
  assign w678[44] = |(datain[135:132] ^ 0);
  assign w678[45] = |(datain[131:128] ^ 0);
  assign w678[46] = |(datain[127:124] ^ 0);
  assign w678[47] = |(datain[123:120] ^ 1);
  assign w678[48] = |(datain[119:116] ^ 12);
  assign w678[49] = |(datain[115:112] ^ 13);
  assign w678[50] = |(datain[111:108] ^ 2);
  assign w678[51] = |(datain[107:104] ^ 1);
  assign w678[52] = |(datain[103:100] ^ 5);
  assign w678[53] = |(datain[99:96] ^ 9);
  assign w678[54] = |(datain[95:92] ^ 5);
  assign w678[55] = |(datain[91:88] ^ 10);
  assign comp[678] = ~(|w678);
  wire [62-1:0] w679;
  assign w679[0] = |(datain[311:308] ^ 0);
  assign w679[1] = |(datain[307:304] ^ 1);
  assign w679[2] = |(datain[303:300] ^ 11);
  assign w679[3] = |(datain[299:296] ^ 8);
  assign w679[4] = |(datain[295:292] ^ 11);
  assign w679[5] = |(datain[291:288] ^ 4);
  assign w679[6] = |(datain[287:284] ^ 4);
  assign w679[7] = |(datain[283:280] ^ 0);
  assign w679[8] = |(datain[279:276] ^ 11);
  assign w679[9] = |(datain[275:272] ^ 9);
  assign w679[10] = |(datain[271:268] ^ 1);
  assign w679[11] = |(datain[267:264] ^ 0);
  assign w679[12] = |(datain[263:260] ^ 0);
  assign w679[13] = |(datain[259:256] ^ 3);
  assign w679[14] = |(datain[255:252] ^ 11);
  assign w679[15] = |(datain[251:248] ^ 10);
  assign w679[16] = |(datain[247:244] ^ 0);
  assign w679[17] = |(datain[243:240] ^ 0);
  assign w679[18] = |(datain[239:236] ^ 0);
  assign w679[19] = |(datain[235:232] ^ 1);
  assign w679[20] = |(datain[231:228] ^ 12);
  assign w679[21] = |(datain[227:224] ^ 13);
  assign w679[22] = |(datain[223:220] ^ 2);
  assign w679[23] = |(datain[219:216] ^ 1);
  assign w679[24] = |(datain[215:212] ^ 11);
  assign w679[25] = |(datain[211:208] ^ 8);
  assign w679[26] = |(datain[207:204] ^ 0);
  assign w679[27] = |(datain[203:200] ^ 0);
  assign w679[28] = |(datain[199:196] ^ 4);
  assign w679[29] = |(datain[195:192] ^ 2);
  assign w679[30] = |(datain[191:188] ^ 3);
  assign w679[31] = |(datain[187:184] ^ 3);
  assign w679[32] = |(datain[183:180] ^ 12);
  assign w679[33] = |(datain[179:176] ^ 9);
  assign w679[34] = |(datain[175:172] ^ 3);
  assign w679[35] = |(datain[171:168] ^ 3);
  assign w679[36] = |(datain[167:164] ^ 13);
  assign w679[37] = |(datain[163:160] ^ 2);
  assign w679[38] = |(datain[159:156] ^ 12);
  assign w679[39] = |(datain[155:152] ^ 13);
  assign w679[40] = |(datain[151:148] ^ 2);
  assign w679[41] = |(datain[147:144] ^ 1);
  assign w679[42] = |(datain[143:140] ^ 11);
  assign w679[43] = |(datain[139:136] ^ 9);
  assign w679[44] = |(datain[135:132] ^ 0);
  assign w679[45] = |(datain[131:128] ^ 3);
  assign w679[46] = |(datain[127:124] ^ 0);
  assign w679[47] = |(datain[123:120] ^ 0);
  assign w679[48] = |(datain[119:116] ^ 11);
  assign w679[49] = |(datain[115:112] ^ 10);
  assign w679[50] = |(datain[111:108] ^ 0);
  assign w679[51] = |(datain[107:104] ^ 0);
  assign w679[52] = |(datain[103:100] ^ 0);
  assign w679[53] = |(datain[99:96] ^ 1);
  assign w679[54] = |(datain[95:92] ^ 11);
  assign w679[55] = |(datain[91:88] ^ 4);
  assign w679[56] = |(datain[87:84] ^ 4);
  assign w679[57] = |(datain[83:80] ^ 0);
  assign w679[58] = |(datain[79:76] ^ 12);
  assign w679[59] = |(datain[75:72] ^ 13);
  assign w679[60] = |(datain[71:68] ^ 2);
  assign w679[61] = |(datain[67:64] ^ 1);
  assign comp[679] = ~(|w679);
  wire [44-1:0] w680;
  assign w680[0] = |(datain[311:308] ^ 11);
  assign w680[1] = |(datain[307:304] ^ 9);
  assign w680[2] = |(datain[303:300] ^ 11);
  assign w680[3] = |(datain[299:296] ^ 11);
  assign w680[4] = |(datain[295:292] ^ 0);
  assign w680[5] = |(datain[291:288] ^ 1);
  assign w680[6] = |(datain[287:284] ^ 11);
  assign w680[7] = |(datain[283:280] ^ 10);
  assign w680[8] = |(datain[279:276] ^ 0);
  assign w680[9] = |(datain[275:272] ^ 0);
  assign w680[10] = |(datain[271:268] ^ 0);
  assign w680[11] = |(datain[267:264] ^ 1);
  assign w680[12] = |(datain[263:260] ^ 12);
  assign w680[13] = |(datain[259:256] ^ 13);
  assign w680[14] = |(datain[255:252] ^ 2);
  assign w680[15] = |(datain[251:248] ^ 1);
  assign w680[16] = |(datain[247:244] ^ 11);
  assign w680[17] = |(datain[243:240] ^ 8);
  assign w680[18] = |(datain[239:236] ^ 0);
  assign w680[19] = |(datain[235:232] ^ 0);
  assign w680[20] = |(datain[231:228] ^ 4);
  assign w680[21] = |(datain[227:224] ^ 2);
  assign w680[22] = |(datain[223:220] ^ 3);
  assign w680[23] = |(datain[219:216] ^ 3);
  assign w680[24] = |(datain[215:212] ^ 12);
  assign w680[25] = |(datain[211:208] ^ 9);
  assign w680[26] = |(datain[207:204] ^ 3);
  assign w680[27] = |(datain[203:200] ^ 3);
  assign w680[28] = |(datain[199:196] ^ 13);
  assign w680[29] = |(datain[195:192] ^ 2);
  assign w680[30] = |(datain[191:188] ^ 12);
  assign w680[31] = |(datain[187:184] ^ 13);
  assign w680[32] = |(datain[183:180] ^ 2);
  assign w680[33] = |(datain[179:176] ^ 1);
  assign w680[34] = |(datain[175:172] ^ 11);
  assign w680[35] = |(datain[171:168] ^ 4);
  assign w680[36] = |(datain[167:164] ^ 4);
  assign w680[37] = |(datain[163:160] ^ 0);
  assign w680[38] = |(datain[159:156] ^ 11);
  assign w680[39] = |(datain[155:152] ^ 9);
  assign w680[40] = |(datain[151:148] ^ 0);
  assign w680[41] = |(datain[147:144] ^ 4);
  assign w680[42] = |(datain[143:140] ^ 0);
  assign w680[43] = |(datain[139:136] ^ 0);
  assign comp[680] = ~(|w680);
  wire [42-1:0] w681;
  assign w681[0] = |(datain[311:308] ^ 2);
  assign w681[1] = |(datain[307:304] ^ 12);
  assign w681[2] = |(datain[303:300] ^ 0);
  assign w681[3] = |(datain[299:296] ^ 4);
  assign w681[4] = |(datain[295:292] ^ 11);
  assign w681[5] = |(datain[291:288] ^ 10);
  assign w681[6] = |(datain[287:284] ^ 0);
  assign w681[7] = |(datain[283:280] ^ 0);
  assign w681[8] = |(datain[279:276] ^ 0);
  assign w681[9] = |(datain[275:272] ^ 1);
  assign w681[10] = |(datain[271:268] ^ 12);
  assign w681[11] = |(datain[267:264] ^ 13);
  assign w681[12] = |(datain[263:260] ^ 2);
  assign w681[13] = |(datain[259:256] ^ 1);
  assign w681[14] = |(datain[255:252] ^ 11);
  assign w681[15] = |(datain[251:248] ^ 8);
  assign w681[16] = |(datain[247:244] ^ 0);
  assign w681[17] = |(datain[243:240] ^ 0);
  assign w681[18] = |(datain[239:236] ^ 4);
  assign w681[19] = |(datain[235:232] ^ 2);
  assign w681[20] = |(datain[231:228] ^ 3);
  assign w681[21] = |(datain[227:224] ^ 3);
  assign w681[22] = |(datain[223:220] ^ 12);
  assign w681[23] = |(datain[219:216] ^ 9);
  assign w681[24] = |(datain[215:212] ^ 3);
  assign w681[25] = |(datain[211:208] ^ 3);
  assign w681[26] = |(datain[207:204] ^ 13);
  assign w681[27] = |(datain[203:200] ^ 2);
  assign w681[28] = |(datain[199:196] ^ 12);
  assign w681[29] = |(datain[195:192] ^ 13);
  assign w681[30] = |(datain[191:188] ^ 2);
  assign w681[31] = |(datain[187:184] ^ 1);
  assign w681[32] = |(datain[183:180] ^ 11);
  assign w681[33] = |(datain[179:176] ^ 4);
  assign w681[34] = |(datain[175:172] ^ 4);
  assign w681[35] = |(datain[171:168] ^ 0);
  assign w681[36] = |(datain[167:164] ^ 11);
  assign w681[37] = |(datain[163:160] ^ 9);
  assign w681[38] = |(datain[159:156] ^ 0);
  assign w681[39] = |(datain[155:152] ^ 4);
  assign w681[40] = |(datain[151:148] ^ 0);
  assign w681[41] = |(datain[147:144] ^ 0);
  assign comp[681] = ~(|w681);
  wire [66-1:0] w682;
  assign w682[0] = |(datain[311:308] ^ 12);
  assign w682[1] = |(datain[307:304] ^ 13);
  assign w682[2] = |(datain[303:300] ^ 2);
  assign w682[3] = |(datain[299:296] ^ 1);
  assign w682[4] = |(datain[295:292] ^ 11);
  assign w682[5] = |(datain[291:288] ^ 8);
  assign w682[6] = |(datain[287:284] ^ 0);
  assign w682[7] = |(datain[283:280] ^ 1);
  assign w682[8] = |(datain[279:276] ^ 5);
  assign w682[9] = |(datain[275:272] ^ 7);
  assign w682[10] = |(datain[271:268] ^ 5);
  assign w682[11] = |(datain[267:264] ^ 10);
  assign w682[12] = |(datain[263:260] ^ 5);
  assign w682[13] = |(datain[259:256] ^ 9);
  assign w682[14] = |(datain[255:252] ^ 12);
  assign w682[15] = |(datain[251:248] ^ 13);
  assign w682[16] = |(datain[247:244] ^ 2);
  assign w682[17] = |(datain[243:240] ^ 1);
  assign w682[18] = |(datain[239:236] ^ 11);
  assign w682[19] = |(datain[235:232] ^ 4);
  assign w682[20] = |(datain[231:228] ^ 3);
  assign w682[21] = |(datain[227:224] ^ 14);
  assign w682[22] = |(datain[223:220] ^ 12);
  assign w682[23] = |(datain[219:216] ^ 13);
  assign w682[24] = |(datain[215:212] ^ 2);
  assign w682[25] = |(datain[211:208] ^ 1);
  assign w682[26] = |(datain[207:204] ^ 2);
  assign w682[27] = |(datain[203:200] ^ 14);
  assign w682[28] = |(datain[199:196] ^ 8);
  assign w682[29] = |(datain[195:192] ^ 0);
  assign w682[30] = |(datain[191:188] ^ 3);
  assign w682[31] = |(datain[187:184] ^ 14);
  assign w682[32] = |(datain[183:180] ^ 0);
  assign w682[33] = |(datain[179:176] ^ 7);
  assign w682[34] = |(datain[175:172] ^ 0);
  assign w682[35] = |(datain[171:168] ^ 1);
  assign w682[36] = |(datain[167:164] ^ 0);
  assign w682[37] = |(datain[163:160] ^ 3);
  assign w682[38] = |(datain[159:156] ^ 7);
  assign w682[39] = |(datain[155:152] ^ 5);
  assign w682[40] = |(datain[151:148] ^ 1);
  assign w682[41] = |(datain[147:144] ^ 12);
  assign w682[42] = |(datain[143:140] ^ 11);
  assign w682[43] = |(datain[139:136] ^ 4);
  assign w682[44] = |(datain[135:132] ^ 1);
  assign w682[45] = |(datain[131:128] ^ 9);
  assign w682[46] = |(datain[127:124] ^ 12);
  assign w682[47] = |(datain[123:120] ^ 13);
  assign w682[48] = |(datain[119:116] ^ 2);
  assign w682[49] = |(datain[115:112] ^ 1);
  assign w682[50] = |(datain[111:108] ^ 11);
  assign w682[51] = |(datain[107:104] ^ 9);
  assign w682[52] = |(datain[103:100] ^ 3);
  assign w682[53] = |(datain[99:96] ^ 3);
  assign w682[54] = |(datain[95:92] ^ 0);
  assign w682[55] = |(datain[91:88] ^ 0);
  assign w682[56] = |(datain[87:84] ^ 11);
  assign w682[57] = |(datain[83:80] ^ 10);
  assign w682[58] = |(datain[79:76] ^ 0);
  assign w682[59] = |(datain[75:72] ^ 0);
  assign w682[60] = |(datain[71:68] ^ 0);
  assign w682[61] = |(datain[67:64] ^ 0);
  assign w682[62] = |(datain[63:60] ^ 12);
  assign w682[63] = |(datain[59:56] ^ 13);
  assign w682[64] = |(datain[55:52] ^ 2);
  assign w682[65] = |(datain[51:48] ^ 6);
  assign comp[682] = ~(|w682);
  wire [44-1:0] w683;
  assign w683[0] = |(datain[311:308] ^ 11);
  assign w683[1] = |(datain[307:304] ^ 9);
  assign w683[2] = |(datain[303:300] ^ 0);
  assign w683[3] = |(datain[299:296] ^ 0);
  assign w683[4] = |(datain[295:292] ^ 0);
  assign w683[5] = |(datain[291:288] ^ 4);
  assign w683[6] = |(datain[287:284] ^ 11);
  assign w683[7] = |(datain[283:280] ^ 10);
  assign w683[8] = |(datain[279:276] ^ 0);
  assign w683[9] = |(datain[275:272] ^ 0);
  assign w683[10] = |(datain[271:268] ^ 0);
  assign w683[11] = |(datain[267:264] ^ 1);
  assign w683[12] = |(datain[263:260] ^ 12);
  assign w683[13] = |(datain[259:256] ^ 13);
  assign w683[14] = |(datain[255:252] ^ 2);
  assign w683[15] = |(datain[251:248] ^ 1);
  assign w683[16] = |(datain[247:244] ^ 11);
  assign w683[17] = |(datain[243:240] ^ 8);
  assign w683[18] = |(datain[239:236] ^ 0);
  assign w683[19] = |(datain[235:232] ^ 0);
  assign w683[20] = |(datain[231:228] ^ 4);
  assign w683[21] = |(datain[227:224] ^ 2);
  assign w683[22] = |(datain[223:220] ^ 3);
  assign w683[23] = |(datain[219:216] ^ 3);
  assign w683[24] = |(datain[215:212] ^ 12);
  assign w683[25] = |(datain[211:208] ^ 9);
  assign w683[26] = |(datain[207:204] ^ 3);
  assign w683[27] = |(datain[203:200] ^ 3);
  assign w683[28] = |(datain[199:196] ^ 13);
  assign w683[29] = |(datain[195:192] ^ 2);
  assign w683[30] = |(datain[191:188] ^ 12);
  assign w683[31] = |(datain[187:184] ^ 13);
  assign w683[32] = |(datain[183:180] ^ 2);
  assign w683[33] = |(datain[179:176] ^ 1);
  assign w683[34] = |(datain[175:172] ^ 11);
  assign w683[35] = |(datain[171:168] ^ 4);
  assign w683[36] = |(datain[167:164] ^ 4);
  assign w683[37] = |(datain[163:160] ^ 0);
  assign w683[38] = |(datain[159:156] ^ 11);
  assign w683[39] = |(datain[155:152] ^ 9);
  assign w683[40] = |(datain[151:148] ^ 0);
  assign w683[41] = |(datain[147:144] ^ 4);
  assign w683[42] = |(datain[143:140] ^ 0);
  assign w683[43] = |(datain[139:136] ^ 0);
  assign comp[683] = ~(|w683);
  wire [42-1:0] w684;
  assign w684[0] = |(datain[311:308] ^ 2);
  assign w684[1] = |(datain[307:304] ^ 2);
  assign w684[2] = |(datain[303:300] ^ 0);
  assign w684[3] = |(datain[299:296] ^ 1);
  assign w684[4] = |(datain[295:292] ^ 11);
  assign w684[5] = |(datain[291:288] ^ 10);
  assign w684[6] = |(datain[287:284] ^ 0);
  assign w684[7] = |(datain[283:280] ^ 0);
  assign w684[8] = |(datain[279:276] ^ 0);
  assign w684[9] = |(datain[275:272] ^ 1);
  assign w684[10] = |(datain[271:268] ^ 12);
  assign w684[11] = |(datain[267:264] ^ 13);
  assign w684[12] = |(datain[263:260] ^ 2);
  assign w684[13] = |(datain[259:256] ^ 1);
  assign w684[14] = |(datain[255:252] ^ 11);
  assign w684[15] = |(datain[251:248] ^ 8);
  assign w684[16] = |(datain[247:244] ^ 0);
  assign w684[17] = |(datain[243:240] ^ 0);
  assign w684[18] = |(datain[239:236] ^ 4);
  assign w684[19] = |(datain[235:232] ^ 2);
  assign w684[20] = |(datain[231:228] ^ 3);
  assign w684[21] = |(datain[227:224] ^ 3);
  assign w684[22] = |(datain[223:220] ^ 12);
  assign w684[23] = |(datain[219:216] ^ 9);
  assign w684[24] = |(datain[215:212] ^ 3);
  assign w684[25] = |(datain[211:208] ^ 3);
  assign w684[26] = |(datain[207:204] ^ 13);
  assign w684[27] = |(datain[203:200] ^ 2);
  assign w684[28] = |(datain[199:196] ^ 12);
  assign w684[29] = |(datain[195:192] ^ 13);
  assign w684[30] = |(datain[191:188] ^ 2);
  assign w684[31] = |(datain[187:184] ^ 1);
  assign w684[32] = |(datain[183:180] ^ 11);
  assign w684[33] = |(datain[179:176] ^ 4);
  assign w684[34] = |(datain[175:172] ^ 4);
  assign w684[35] = |(datain[171:168] ^ 0);
  assign w684[36] = |(datain[167:164] ^ 11);
  assign w684[37] = |(datain[163:160] ^ 9);
  assign w684[38] = |(datain[159:156] ^ 0);
  assign w684[39] = |(datain[155:152] ^ 4);
  assign w684[40] = |(datain[151:148] ^ 0);
  assign w684[41] = |(datain[147:144] ^ 0);
  assign comp[684] = ~(|w684);
  wire [44-1:0] w685;
  assign w685[0] = |(datain[311:308] ^ 3);
  assign w685[1] = |(datain[307:304] ^ 3);
  assign w685[2] = |(datain[303:300] ^ 12);
  assign w685[3] = |(datain[299:296] ^ 9);
  assign w685[4] = |(datain[295:292] ^ 12);
  assign w685[5] = |(datain[291:288] ^ 13);
  assign w685[6] = |(datain[287:284] ^ 2);
  assign w685[7] = |(datain[283:280] ^ 1);
  assign w685[8] = |(datain[279:276] ^ 8);
  assign w685[9] = |(datain[275:272] ^ 11);
  assign w685[10] = |(datain[271:268] ^ 13);
  assign w685[11] = |(datain[267:264] ^ 8);
  assign w685[12] = |(datain[263:260] ^ 11);
  assign w685[13] = |(datain[259:256] ^ 4);
  assign w685[14] = |(datain[255:252] ^ 4);
  assign w685[15] = |(datain[251:248] ^ 0);
  assign w685[16] = |(datain[247:244] ^ 11);
  assign w685[17] = |(datain[243:240] ^ 9);
  assign w685[18] = |(datain[239:236] ^ 0);
  assign w685[19] = |(datain[235:232] ^ 7);
  assign w685[20] = |(datain[231:228] ^ 0);
  assign w685[21] = |(datain[227:224] ^ 14);
  assign w685[22] = |(datain[223:220] ^ 8);
  assign w685[23] = |(datain[219:216] ^ 13);
  assign w685[24] = |(datain[215:212] ^ 9);
  assign w685[25] = |(datain[211:208] ^ 6);
  assign w685[26] = |(datain[207:204] ^ 3);
  assign w685[27] = |(datain[203:200] ^ 1);
  assign w685[28] = |(datain[199:196] ^ 0);
  assign w685[29] = |(datain[195:192] ^ 2);
  assign w685[30] = |(datain[191:188] ^ 12);
  assign w685[31] = |(datain[187:184] ^ 13);
  assign w685[32] = |(datain[183:180] ^ 2);
  assign w685[33] = |(datain[179:176] ^ 1);
  assign w685[34] = |(datain[175:172] ^ 11);
  assign w685[35] = |(datain[171:168] ^ 4);
  assign w685[36] = |(datain[167:164] ^ 3);
  assign w685[37] = |(datain[163:160] ^ 14);
  assign w685[38] = |(datain[159:156] ^ 12);
  assign w685[39] = |(datain[155:152] ^ 13);
  assign w685[40] = |(datain[151:148] ^ 2);
  assign w685[41] = |(datain[147:144] ^ 1);
  assign w685[42] = |(datain[143:140] ^ 12);
  assign w685[43] = |(datain[139:136] ^ 3);
  assign comp[685] = ~(|w685);
  wire [46-1:0] w686;
  assign w686[0] = |(datain[311:308] ^ 15);
  assign w686[1] = |(datain[307:304] ^ 15);
  assign w686[2] = |(datain[303:300] ^ 11);
  assign w686[3] = |(datain[299:296] ^ 10);
  assign w686[4] = |(datain[295:292] ^ 8);
  assign w686[5] = |(datain[291:288] ^ 0);
  assign w686[6] = |(datain[287:284] ^ 0);
  assign w686[7] = |(datain[283:280] ^ 0);
  assign w686[8] = |(datain[279:276] ^ 11);
  assign w686[9] = |(datain[275:272] ^ 11);
  assign w686[10] = |(datain[271:268] ^ 0);
  assign w686[11] = |(datain[267:264] ^ 0);
  assign w686[12] = |(datain[263:260] ^ 0);
  assign w686[13] = |(datain[259:256] ^ 7);
  assign w686[14] = |(datain[255:252] ^ 8);
  assign w686[15] = |(datain[251:248] ^ 11);
  assign w686[16] = |(datain[247:244] ^ 12);
  assign w686[17] = |(datain[243:240] ^ 15);
  assign w686[18] = |(datain[239:236] ^ 8);
  assign w686[19] = |(datain[235:232] ^ 3);
  assign w686[20] = |(datain[231:228] ^ 12);
  assign w686[21] = |(datain[227:224] ^ 1);
  assign w686[22] = |(datain[223:220] ^ 0);
  assign w686[23] = |(datain[219:216] ^ 3);
  assign w686[24] = |(datain[215:212] ^ 11);
  assign w686[25] = |(datain[211:208] ^ 8);
  assign w686[26] = |(datain[207:204] ^ 0);
  assign w686[27] = |(datain[203:200] ^ 1);
  assign w686[28] = |(datain[199:196] ^ 0);
  assign w686[29] = |(datain[195:192] ^ 2);
  assign w686[30] = |(datain[191:188] ^ 12);
  assign w686[31] = |(datain[187:184] ^ 13);
  assign w686[32] = |(datain[183:180] ^ 1);
  assign w686[33] = |(datain[179:176] ^ 3);
  assign w686[34] = |(datain[175:172] ^ 8);
  assign w686[35] = |(datain[171:168] ^ 1);
  assign w686[36] = |(datain[167:164] ^ 14);
  assign w686[37] = |(datain[163:160] ^ 11);
  assign w686[38] = |(datain[159:156] ^ 0);
  assign w686[39] = |(datain[155:152] ^ 0);
  assign w686[40] = |(datain[151:148] ^ 0);
  assign w686[41] = |(datain[147:144] ^ 2);
  assign w686[42] = |(datain[143:140] ^ 4);
  assign w686[43] = |(datain[139:136] ^ 7);
  assign w686[44] = |(datain[135:132] ^ 8);
  assign w686[45] = |(datain[131:128] ^ 3);
  assign comp[686] = ~(|w686);
  wire [74-1:0] w687;
  assign w687[0] = |(datain[311:308] ^ 0);
  assign w687[1] = |(datain[307:304] ^ 2);
  assign w687[2] = |(datain[303:300] ^ 10);
  assign w687[3] = |(datain[299:296] ^ 1);
  assign w687[4] = |(datain[295:292] ^ 0);
  assign w687[5] = |(datain[291:288] ^ 13);
  assign w687[6] = |(datain[287:284] ^ 0);
  assign w687[7] = |(datain[283:280] ^ 2);
  assign w687[8] = |(datain[279:276] ^ 2);
  assign w687[9] = |(datain[275:272] ^ 11);
  assign w687[10] = |(datain[271:268] ^ 0);
  assign w687[11] = |(datain[267:264] ^ 6);
  assign w687[12] = |(datain[263:260] ^ 0);
  assign w687[13] = |(datain[259:256] ^ 1);
  assign w687[14] = |(datain[255:252] ^ 0);
  assign w687[15] = |(datain[251:248] ^ 2);
  assign w687[16] = |(datain[247:244] ^ 10);
  assign w687[17] = |(datain[243:240] ^ 3);
  assign w687[18] = |(datain[239:236] ^ 3);
  assign w687[19] = |(datain[235:232] ^ 0);
  assign w687[20] = |(datain[231:228] ^ 0);
  assign w687[21] = |(datain[227:224] ^ 0);
  assign w687[22] = |(datain[223:220] ^ 10);
  assign w687[23] = |(datain[219:216] ^ 1);
  assign w687[24] = |(datain[215:212] ^ 15);
  assign w687[25] = |(datain[211:208] ^ 15);
  assign w687[26] = |(datain[207:204] ^ 0);
  assign w687[27] = |(datain[203:200] ^ 1);
  assign w687[28] = |(datain[199:196] ^ 10);
  assign w687[29] = |(datain[195:192] ^ 3);
  assign w687[30] = |(datain[191:188] ^ 2);
  assign w687[31] = |(datain[187:184] ^ 12);
  assign w687[32] = |(datain[183:180] ^ 0);
  assign w687[33] = |(datain[179:176] ^ 0);
  assign w687[34] = |(datain[175:172] ^ 11);
  assign w687[35] = |(datain[171:168] ^ 4);
  assign w687[36] = |(datain[167:164] ^ 4);
  assign w687[37] = |(datain[163:160] ^ 0);
  assign w687[38] = |(datain[159:156] ^ 8);
  assign w687[39] = |(datain[155:152] ^ 11);
  assign w687[40] = |(datain[151:148] ^ 1);
  assign w687[41] = |(datain[147:144] ^ 14);
  assign w687[42] = |(datain[143:140] ^ 14);
  assign w687[43] = |(datain[139:136] ^ 9);
  assign w687[44] = |(datain[135:132] ^ 0);
  assign w687[45] = |(datain[131:128] ^ 1);
  assign w687[46] = |(datain[127:124] ^ 11);
  assign w687[47] = |(datain[123:120] ^ 9);
  assign w687[48] = |(datain[119:116] ^ 2);
  assign w687[49] = |(datain[115:112] ^ 6);
  assign w687[50] = |(datain[111:108] ^ 0);
  assign w687[51] = |(datain[107:104] ^ 2);
  assign w687[52] = |(datain[103:100] ^ 11);
  assign w687[53] = |(datain[99:96] ^ 10);
  assign w687[54] = |(datain[95:92] ^ 0);
  assign w687[55] = |(datain[91:88] ^ 0);
  assign w687[56] = |(datain[87:84] ^ 0);
  assign w687[57] = |(datain[83:80] ^ 0);
  assign w687[58] = |(datain[79:76] ^ 12);
  assign w687[59] = |(datain[75:72] ^ 13);
  assign w687[60] = |(datain[71:68] ^ 2);
  assign w687[61] = |(datain[67:64] ^ 1);
  assign w687[62] = |(datain[63:60] ^ 7);
  assign w687[63] = |(datain[59:56] ^ 3);
  assign w687[64] = |(datain[55:52] ^ 0);
  assign w687[65] = |(datain[51:48] ^ 3);
  assign w687[66] = |(datain[47:44] ^ 14);
  assign w687[67] = |(datain[43:40] ^ 11);
  assign w687[68] = |(datain[39:36] ^ 2);
  assign w687[69] = |(datain[35:32] ^ 13);
  assign w687[70] = |(datain[31:28] ^ 9);
  assign w687[71] = |(datain[27:24] ^ 0);
  assign w687[72] = |(datain[23:20] ^ 11);
  assign w687[73] = |(datain[19:16] ^ 8);
  assign comp[687] = ~(|w687);
  wire [34-1:0] w688;
  assign w688[0] = |(datain[311:308] ^ 0);
  assign w688[1] = |(datain[307:304] ^ 10);
  assign w688[2] = |(datain[303:300] ^ 0);
  assign w688[3] = |(datain[299:296] ^ 0);
  assign w688[4] = |(datain[295:292] ^ 0);
  assign w688[5] = |(datain[291:288] ^ 0);
  assign w688[6] = |(datain[287:284] ^ 11);
  assign w688[7] = |(datain[283:280] ^ 11);
  assign w688[8] = |(datain[279:276] ^ 1);
  assign w688[9] = |(datain[275:272] ^ 14);
  assign w688[10] = |(datain[271:268] ^ 0);
  assign w688[11] = |(datain[267:264] ^ 2);
  assign w688[12] = |(datain[263:260] ^ 14);
  assign w688[13] = |(datain[259:256] ^ 11);
  assign w688[14] = |(datain[255:252] ^ 0);
  assign w688[15] = |(datain[251:248] ^ 7);
  assign w688[16] = |(datain[247:244] ^ 9);
  assign w688[17] = |(datain[243:240] ^ 0);
  assign w688[18] = |(datain[239:236] ^ 14);
  assign w688[19] = |(datain[235:232] ^ 10);
  assign w688[20] = |(datain[231:228] ^ 2);
  assign w688[21] = |(datain[227:224] ^ 14);
  assign w688[22] = |(datain[223:220] ^ 8);
  assign w688[23] = |(datain[219:216] ^ 0);
  assign w688[24] = |(datain[215:212] ^ 3);
  assign w688[25] = |(datain[211:208] ^ 7);
  assign w688[26] = |(datain[207:204] ^ 0);
  assign w688[27] = |(datain[203:200] ^ 0);
  assign w688[28] = |(datain[199:196] ^ 4);
  assign w688[29] = |(datain[195:192] ^ 3);
  assign w688[30] = |(datain[191:188] ^ 14);
  assign w688[31] = |(datain[187:184] ^ 2);
  assign w688[32] = |(datain[183:180] ^ 15);
  assign w688[33] = |(datain[179:176] ^ 9);
  assign comp[688] = ~(|w688);
  wire [44-1:0] w689;
  assign w689[0] = |(datain[311:308] ^ 5);
  assign w689[1] = |(datain[307:304] ^ 14);
  assign w689[2] = |(datain[303:300] ^ 0);
  assign w689[3] = |(datain[299:296] ^ 1);
  assign w689[4] = |(datain[295:292] ^ 8);
  assign w689[5] = |(datain[291:288] ^ 13);
  assign w689[6] = |(datain[287:284] ^ 7);
  assign w689[7] = |(datain[283:280] ^ 4);
  assign w689[8] = |(datain[279:276] ^ 15);
  assign w689[9] = |(datain[275:272] ^ 12);
  assign w689[10] = |(datain[271:268] ^ 11);
  assign w689[11] = |(datain[267:264] ^ 0);
  assign w689[12] = |(datain[263:260] ^ 9);
  assign w689[13] = |(datain[259:256] ^ 4);
  assign w689[14] = |(datain[255:252] ^ 0);
  assign w689[15] = |(datain[251:248] ^ 14);
  assign w689[16] = |(datain[247:244] ^ 1);
  assign w689[17] = |(datain[243:240] ^ 7);
  assign w689[18] = |(datain[239:236] ^ 8);
  assign w689[19] = |(datain[235:232] ^ 13);
  assign w689[20] = |(datain[231:228] ^ 6);
  assign w689[21] = |(datain[227:224] ^ 4);
  assign w689[22] = |(datain[223:220] ^ 2);
  assign w689[23] = |(datain[219:216] ^ 0);
  assign w689[24] = |(datain[215:212] ^ 5);
  assign w689[25] = |(datain[211:208] ^ 10);
  assign w689[26] = |(datain[207:204] ^ 3);
  assign w689[27] = |(datain[203:200] ^ 2);
  assign w689[28] = |(datain[199:196] ^ 15);
  assign w689[29] = |(datain[195:192] ^ 0);
  assign w689[30] = |(datain[191:188] ^ 3);
  assign w689[31] = |(datain[187:184] ^ 2);
  assign w689[32] = |(datain[183:180] ^ 13);
  assign w689[33] = |(datain[179:176] ^ 0);
  assign w689[34] = |(datain[175:172] ^ 5);
  assign w689[35] = |(datain[171:168] ^ 2);
  assign w689[36] = |(datain[167:164] ^ 4);
  assign w689[37] = |(datain[163:160] ^ 4);
  assign w689[38] = |(datain[159:156] ^ 4);
  assign w689[39] = |(datain[155:152] ^ 4);
  assign w689[40] = |(datain[151:148] ^ 14);
  assign w689[41] = |(datain[147:144] ^ 2);
  assign w689[42] = |(datain[143:140] ^ 15);
  assign w689[43] = |(datain[139:136] ^ 6);
  assign comp[689] = ~(|w689);
  wire [44-1:0] w690;
  assign w690[0] = |(datain[311:308] ^ 12);
  assign w690[1] = |(datain[307:304] ^ 13);
  assign w690[2] = |(datain[303:300] ^ 2);
  assign w690[3] = |(datain[299:296] ^ 1);
  assign w690[4] = |(datain[295:292] ^ 8);
  assign w690[5] = |(datain[291:288] ^ 0);
  assign w690[6] = |(datain[287:284] ^ 15);
  assign w690[7] = |(datain[283:280] ^ 12);
  assign w690[8] = |(datain[279:276] ^ 14);
  assign w690[9] = |(datain[275:272] ^ 14);
  assign w690[10] = |(datain[271:268] ^ 7);
  assign w690[11] = |(datain[267:264] ^ 4);
  assign w690[12] = |(datain[263:260] ^ 0);
  assign w690[13] = |(datain[259:256] ^ 6);
  assign w690[14] = |(datain[255:252] ^ 8);
  assign w690[15] = |(datain[251:248] ^ 3);
  assign w690[16] = |(datain[247:244] ^ 14);
  assign w690[17] = |(datain[243:240] ^ 14);
  assign w690[18] = |(datain[239:236] ^ 0);
  assign w690[19] = |(datain[235:232] ^ 6);
  assign w690[20] = |(datain[231:228] ^ 14);
  assign w690[21] = |(datain[227:224] ^ 8);
  assign w690[22] = |(datain[223:220] ^ 0);
  assign w690[23] = |(datain[219:216] ^ 8);
  assign w690[24] = |(datain[215:212] ^ 0);
  assign w690[25] = |(datain[211:208] ^ 0);
  assign w690[26] = |(datain[207:204] ^ 11);
  assign w690[27] = |(datain[203:200] ^ 15);
  assign w690[28] = |(datain[199:196] ^ 0);
  assign w690[29] = |(datain[195:192] ^ 0);
  assign w690[30] = |(datain[191:188] ^ 0);
  assign w690[31] = |(datain[187:184] ^ 1);
  assign w690[32] = |(datain[183:180] ^ 5);
  assign w690[33] = |(datain[179:176] ^ 7);
  assign w690[34] = |(datain[175:172] ^ 12);
  assign w690[35] = |(datain[171:168] ^ 3);
  assign w690[36] = |(datain[167:164] ^ 11);
  assign w690[37] = |(datain[163:160] ^ 0);
  assign w690[38] = |(datain[159:156] ^ 0);
  assign w690[39] = |(datain[155:152] ^ 3);
  assign w690[40] = |(datain[151:148] ^ 12);
  assign w690[41] = |(datain[147:144] ^ 15);
  assign w690[42] = |(datain[143:140] ^ 0);
  assign w690[43] = |(datain[139:136] ^ 6);
  assign comp[690] = ~(|w690);
  wire [74-1:0] w691;
  assign w691[0] = |(datain[311:308] ^ 11);
  assign w691[1] = |(datain[307:304] ^ 6);
  assign w691[2] = |(datain[303:300] ^ 0);
  assign w691[3] = |(datain[299:296] ^ 9);
  assign w691[4] = |(datain[295:292] ^ 0);
  assign w691[5] = |(datain[291:288] ^ 1);
  assign w691[6] = |(datain[287:284] ^ 11);
  assign w691[7] = |(datain[283:280] ^ 15);
  assign w691[8] = |(datain[279:276] ^ 11);
  assign w691[9] = |(datain[275:272] ^ 14);
  assign w691[10] = |(datain[271:268] ^ 15);
  assign w691[11] = |(datain[267:264] ^ 9);
  assign w691[12] = |(datain[263:260] ^ 11);
  assign w691[13] = |(datain[259:256] ^ 9);
  assign w691[14] = |(datain[255:252] ^ 0);
  assign w691[15] = |(datain[251:248] ^ 11);
  assign w691[16] = |(datain[247:244] ^ 0);
  assign w691[17] = |(datain[243:240] ^ 1);
  assign w691[18] = |(datain[239:236] ^ 15);
  assign w691[19] = |(datain[235:232] ^ 3);
  assign w691[20] = |(datain[231:228] ^ 10);
  assign w691[21] = |(datain[227:224] ^ 4);
  assign w691[22] = |(datain[223:220] ^ 11);
  assign w691[23] = |(datain[219:216] ^ 14);
  assign w691[24] = |(datain[215:212] ^ 14);
  assign w691[25] = |(datain[211:208] ^ 2);
  assign w691[26] = |(datain[207:204] ^ 15);
  assign w691[27] = |(datain[203:200] ^ 9);
  assign w691[28] = |(datain[199:196] ^ 14);
  assign w691[29] = |(datain[195:192] ^ 8);
  assign w691[30] = |(datain[191:188] ^ 5);
  assign w691[31] = |(datain[187:184] ^ 11);
  assign w691[32] = |(datain[183:180] ^ 15);
  assign w691[33] = |(datain[179:176] ^ 15);
  assign w691[34] = |(datain[175:172] ^ 11);
  assign w691[35] = |(datain[171:168] ^ 4);
  assign w691[36] = |(datain[167:164] ^ 4);
  assign w691[37] = |(datain[163:160] ^ 0);
  assign w691[38] = |(datain[159:156] ^ 11);
  assign w691[39] = |(datain[155:152] ^ 10);
  assign w691[40] = |(datain[151:148] ^ 11);
  assign w691[41] = |(datain[147:144] ^ 14);
  assign w691[42] = |(datain[143:140] ^ 15);
  assign w691[43] = |(datain[139:136] ^ 9);
  assign w691[44] = |(datain[135:132] ^ 11);
  assign w691[45] = |(datain[131:128] ^ 9);
  assign w691[46] = |(datain[127:124] ^ 0);
  assign w691[47] = |(datain[123:120] ^ 11);
  assign w691[48] = |(datain[119:116] ^ 0);
  assign w691[49] = |(datain[115:112] ^ 1);
  assign w691[50] = |(datain[111:108] ^ 12);
  assign w691[51] = |(datain[107:104] ^ 13);
  assign w691[52] = |(datain[103:100] ^ 2);
  assign w691[53] = |(datain[99:96] ^ 1);
  assign w691[54] = |(datain[95:92] ^ 11);
  assign w691[55] = |(datain[91:88] ^ 8);
  assign w691[56] = |(datain[87:84] ^ 0);
  assign w691[57] = |(datain[83:80] ^ 0);
  assign w691[58] = |(datain[79:76] ^ 4);
  assign w691[59] = |(datain[75:72] ^ 2);
  assign w691[60] = |(datain[71:68] ^ 14);
  assign w691[61] = |(datain[67:64] ^ 8);
  assign w691[62] = |(datain[63:60] ^ 1);
  assign w691[63] = |(datain[59:56] ^ 12);
  assign w691[64] = |(datain[55:52] ^ 0);
  assign w691[65] = |(datain[51:48] ^ 0);
  assign w691[66] = |(datain[47:44] ^ 11);
  assign w691[67] = |(datain[43:40] ^ 4);
  assign w691[68] = |(datain[39:36] ^ 4);
  assign w691[69] = |(datain[35:32] ^ 0);
  assign w691[70] = |(datain[31:28] ^ 11);
  assign w691[71] = |(datain[27:24] ^ 9);
  assign w691[72] = |(datain[23:20] ^ 0);
  assign w691[73] = |(datain[19:16] ^ 3);
  assign comp[691] = ~(|w691);
  wire [66-1:0] w692;
  assign w692[0] = |(datain[311:308] ^ 5);
  assign w692[1] = |(datain[307:304] ^ 11);
  assign w692[2] = |(datain[303:300] ^ 8);
  assign w692[3] = |(datain[299:296] ^ 1);
  assign w692[4] = |(datain[295:292] ^ 14);
  assign w692[5] = |(datain[291:288] ^ 11);
  assign w692[6] = |(datain[287:284] ^ 1);
  assign w692[7] = |(datain[283:280] ^ 2);
  assign w692[8] = |(datain[279:276] ^ 0);
  assign w692[9] = |(datain[275:272] ^ 1);
  assign w692[10] = |(datain[271:268] ^ 8);
  assign w692[11] = |(datain[267:264] ^ 11);
  assign w692[12] = |(datain[263:260] ^ 14);
  assign w692[13] = |(datain[259:256] ^ 11);
  assign w692[14] = |(datain[255:252] ^ 8);
  assign w692[15] = |(datain[251:248] ^ 13);
  assign w692[16] = |(datain[247:244] ^ 11);
  assign w692[17] = |(datain[243:240] ^ 6);
  assign w692[18] = |(datain[239:236] ^ 3);
  assign w692[19] = |(datain[235:232] ^ 3);
  assign w692[20] = |(datain[231:228] ^ 0);
  assign w692[21] = |(datain[227:224] ^ 1);
  assign w692[22] = |(datain[223:220] ^ 5);
  assign w692[23] = |(datain[219:216] ^ 6);
  assign w692[24] = |(datain[215:212] ^ 8);
  assign w692[25] = |(datain[211:208] ^ 11);
  assign w692[26] = |(datain[207:204] ^ 9);
  assign w692[27] = |(datain[203:200] ^ 6);
  assign w692[28] = |(datain[199:196] ^ 2);
  assign w692[29] = |(datain[195:192] ^ 13);
  assign w692[30] = |(datain[191:188] ^ 0);
  assign w692[31] = |(datain[187:184] ^ 2);
  assign w692[32] = |(datain[183:180] ^ 11);
  assign w692[33] = |(datain[179:176] ^ 9);
  assign w692[34] = |(datain[175:172] ^ 7);
  assign w692[35] = |(datain[171:168] ^ 10);
  assign w692[36] = |(datain[167:164] ^ 0);
  assign w692[37] = |(datain[163:160] ^ 0);
  assign w692[38] = |(datain[159:156] ^ 8);
  assign w692[39] = |(datain[155:152] ^ 11);
  assign w692[40] = |(datain[151:148] ^ 15);
  assign w692[41] = |(datain[147:144] ^ 14);
  assign w692[42] = |(datain[143:140] ^ 8);
  assign w692[43] = |(datain[139:136] ^ 4);
  assign w692[44] = |(datain[135:132] ^ 15);
  assign w692[45] = |(datain[131:128] ^ 15);
  assign w692[46] = |(datain[127:124] ^ 15);
  assign w692[47] = |(datain[123:120] ^ 12);
  assign w692[48] = |(datain[119:116] ^ 10);
  assign w692[49] = |(datain[115:112] ^ 13);
  assign w692[50] = |(datain[111:108] ^ 3);
  assign w692[51] = |(datain[107:104] ^ 3);
  assign w692[52] = |(datain[103:100] ^ 12);
  assign w692[53] = |(datain[99:96] ^ 2);
  assign w692[54] = |(datain[95:92] ^ 10);
  assign w692[55] = |(datain[91:88] ^ 11);
  assign w692[56] = |(datain[87:84] ^ 8);
  assign w692[57] = |(datain[83:80] ^ 4);
  assign w692[58] = |(datain[79:76] ^ 13);
  assign w692[59] = |(datain[75:72] ^ 8);
  assign w692[60] = |(datain[71:68] ^ 14);
  assign w692[61] = |(datain[67:64] ^ 2);
  assign w692[62] = |(datain[63:60] ^ 15);
  assign w692[63] = |(datain[59:56] ^ 8);
  assign w692[64] = |(datain[55:52] ^ 12);
  assign w692[65] = |(datain[51:48] ^ 3);
  assign comp[692] = ~(|w692);
  wire [74-1:0] w693;
  assign w693[0] = |(datain[311:308] ^ 5);
  assign w693[1] = |(datain[307:304] ^ 11);
  assign w693[2] = |(datain[303:300] ^ 8);
  assign w693[3] = |(datain[299:296] ^ 1);
  assign w693[4] = |(datain[295:292] ^ 14);
  assign w693[5] = |(datain[291:288] ^ 11);
  assign w693[6] = |(datain[287:284] ^ 0);
  assign w693[7] = |(datain[283:280] ^ 14);
  assign w693[8] = |(datain[279:276] ^ 0);
  assign w693[9] = |(datain[275:272] ^ 0);
  assign w693[10] = |(datain[271:268] ^ 5);
  assign w693[11] = |(datain[267:264] ^ 3);
  assign w693[12] = |(datain[263:260] ^ 3);
  assign w693[13] = |(datain[259:256] ^ 3);
  assign w693[14] = |(datain[255:252] ^ 12);
  assign w693[15] = |(datain[251:248] ^ 0);
  assign w693[16] = |(datain[247:244] ^ 8);
  assign w693[17] = |(datain[243:240] ^ 14);
  assign w693[18] = |(datain[239:236] ^ 13);
  assign w693[19] = |(datain[235:232] ^ 8);
  assign w693[20] = |(datain[231:228] ^ 10);
  assign w693[21] = |(datain[227:224] ^ 1);
  assign w693[22] = |(datain[223:220] ^ 1);
  assign w693[23] = |(datain[219:216] ^ 3);
  assign w693[24] = |(datain[215:212] ^ 0);
  assign w693[25] = |(datain[211:208] ^ 4);
  assign w693[26] = |(datain[207:204] ^ 4);
  assign w693[27] = |(datain[203:200] ^ 8);
  assign w693[28] = |(datain[199:196] ^ 4);
  assign w693[29] = |(datain[195:192] ^ 8);
  assign w693[30] = |(datain[191:188] ^ 10);
  assign w693[31] = |(datain[187:184] ^ 3);
  assign w693[32] = |(datain[183:180] ^ 1);
  assign w693[33] = |(datain[179:176] ^ 3);
  assign w693[34] = |(datain[175:172] ^ 0);
  assign w693[35] = |(datain[171:168] ^ 4);
  assign w693[36] = |(datain[167:164] ^ 11);
  assign w693[37] = |(datain[163:160] ^ 1);
  assign w693[38] = |(datain[159:156] ^ 0);
  assign w693[39] = |(datain[155:152] ^ 6);
  assign w693[40] = |(datain[151:148] ^ 13);
  assign w693[41] = |(datain[147:144] ^ 3);
  assign w693[42] = |(datain[143:140] ^ 14);
  assign w693[43] = |(datain[139:136] ^ 0);
  assign w693[44] = |(datain[135:132] ^ 8);
  assign w693[45] = |(datain[131:128] ^ 14);
  assign w693[46] = |(datain[127:124] ^ 12);
  assign w693[47] = |(datain[123:120] ^ 0);
  assign w693[48] = |(datain[119:116] ^ 3);
  assign w693[49] = |(datain[115:112] ^ 3);
  assign w693[50] = |(datain[111:108] ^ 13);
  assign w693[51] = |(datain[107:104] ^ 11);
  assign w693[52] = |(datain[103:100] ^ 11);
  assign w693[53] = |(datain[99:96] ^ 8);
  assign w693[54] = |(datain[95:92] ^ 0);
  assign w693[55] = |(datain[91:88] ^ 4);
  assign w693[56] = |(datain[87:84] ^ 0);
  assign w693[57] = |(datain[83:80] ^ 2);
  assign w693[58] = |(datain[79:76] ^ 14);
  assign w693[59] = |(datain[75:72] ^ 8);
  assign w693[60] = |(datain[71:68] ^ 9);
  assign w693[61] = |(datain[67:64] ^ 7);
  assign w693[62] = |(datain[63:60] ^ 0);
  assign w693[63] = |(datain[59:56] ^ 0);
  assign w693[64] = |(datain[55:52] ^ 7);
  assign w693[65] = |(datain[51:48] ^ 3);
  assign w693[66] = |(datain[47:44] ^ 0);
  assign w693[67] = |(datain[43:40] ^ 6);
  assign w693[68] = |(datain[39:36] ^ 3);
  assign w693[69] = |(datain[35:32] ^ 3);
  assign w693[70] = |(datain[31:28] ^ 12);
  assign w693[71] = |(datain[27:24] ^ 0);
  assign w693[72] = |(datain[23:20] ^ 12);
  assign w693[73] = |(datain[19:16] ^ 13);
  assign comp[693] = ~(|w693);
  wire [42-1:0] w694;
  assign w694[0] = |(datain[311:308] ^ 0);
  assign w694[1] = |(datain[307:304] ^ 1);
  assign w694[2] = |(datain[303:300] ^ 11);
  assign w694[3] = |(datain[299:296] ^ 14);
  assign w694[4] = |(datain[295:292] ^ 8);
  assign w694[5] = |(datain[291:288] ^ 2);
  assign w694[6] = |(datain[287:284] ^ 0);
  assign w694[7] = |(datain[283:280] ^ 1);
  assign w694[8] = |(datain[279:276] ^ 0);
  assign w694[9] = |(datain[275:272] ^ 3);
  assign w694[10] = |(datain[271:268] ^ 15);
  assign w694[11] = |(datain[267:264] ^ 3);
  assign w694[12] = |(datain[263:260] ^ 11);
  assign w694[13] = |(datain[259:256] ^ 10);
  assign w694[14] = |(datain[255:252] ^ 10);
  assign w694[15] = |(datain[251:248] ^ 15);
  assign w694[16] = |(datain[247:244] ^ 0);
  assign w694[17] = |(datain[243:240] ^ 5);
  assign w694[18] = |(datain[239:236] ^ 0);
  assign w694[19] = |(datain[235:232] ^ 3);
  assign w694[20] = |(datain[231:228] ^ 13);
  assign w694[21] = |(datain[227:224] ^ 3);
  assign w694[22] = |(datain[223:220] ^ 8);
  assign w694[23] = |(datain[219:216] ^ 1);
  assign w694[24] = |(datain[215:212] ^ 3);
  assign w694[25] = |(datain[211:208] ^ 4);
  assign w694[26] = |(datain[207:204] ^ 5);
  assign w694[27] = |(datain[203:200] ^ 0);
  assign w694[28] = |(datain[199:196] ^ 8);
  assign w694[29] = |(datain[195:192] ^ 0);
  assign w694[30] = |(datain[191:188] ^ 4);
  assign w694[31] = |(datain[187:184] ^ 6);
  assign w694[32] = |(datain[183:180] ^ 3);
  assign w694[33] = |(datain[179:176] ^ 11);
  assign w694[34] = |(datain[175:172] ^ 15);
  assign w694[35] = |(datain[171:168] ^ 2);
  assign w694[36] = |(datain[167:164] ^ 7);
  assign w694[37] = |(datain[163:160] ^ 5);
  assign w694[38] = |(datain[159:156] ^ 15);
  assign w694[39] = |(datain[155:152] ^ 7);
  assign w694[40] = |(datain[151:148] ^ 14);
  assign w694[41] = |(datain[147:144] ^ 9);
  assign comp[694] = ~(|w694);
  wire [76-1:0] w695;
  assign w695[0] = |(datain[311:308] ^ 5);
  assign w695[1] = |(datain[307:304] ^ 1);
  assign w695[2] = |(datain[303:300] ^ 0);
  assign w695[3] = |(datain[299:296] ^ 0);
  assign w695[4] = |(datain[295:292] ^ 5);
  assign w695[5] = |(datain[291:288] ^ 13);
  assign w695[6] = |(datain[287:284] ^ 5);
  assign w695[7] = |(datain[283:280] ^ 11);
  assign w695[8] = |(datain[279:276] ^ 8);
  assign w695[9] = |(datain[275:272] ^ 13);
  assign w695[10] = |(datain[271:268] ^ 11);
  assign w695[11] = |(datain[267:264] ^ 6);
  assign w695[12] = |(datain[263:260] ^ 15);
  assign w695[13] = |(datain[259:256] ^ 13);
  assign w695[14] = |(datain[255:252] ^ 15);
  assign w695[15] = |(datain[251:248] ^ 15);
  assign w695[16] = |(datain[247:244] ^ 15);
  assign w695[17] = |(datain[243:240] ^ 12);
  assign w695[18] = |(datain[239:236] ^ 8);
  assign w695[19] = |(datain[235:232] ^ 6);
  assign w695[20] = |(datain[231:228] ^ 12);
  assign w695[21] = |(datain[227:224] ^ 4);
  assign w695[22] = |(datain[223:220] ^ 8);
  assign w695[23] = |(datain[219:216] ^ 7);
  assign w695[24] = |(datain[215:212] ^ 13);
  assign w695[25] = |(datain[211:208] ^ 1);
  assign w695[26] = |(datain[207:204] ^ 5);
  assign w695[27] = |(datain[203:200] ^ 1);
  assign w695[28] = |(datain[199:196] ^ 10);
  assign w695[29] = |(datain[195:192] ^ 12);
  assign w695[30] = |(datain[191:188] ^ 3);
  assign w695[31] = |(datain[187:184] ^ 2);
  assign w695[32] = |(datain[183:180] ^ 12);
  assign w695[33] = |(datain[179:176] ^ 4);
  assign w695[34] = |(datain[175:172] ^ 10);
  assign w695[35] = |(datain[171:168] ^ 10);
  assign w695[36] = |(datain[167:164] ^ 14);
  assign w695[37] = |(datain[163:160] ^ 2);
  assign w695[38] = |(datain[159:156] ^ 15);
  assign w695[39] = |(datain[155:152] ^ 10);
  assign w695[40] = |(datain[151:148] ^ 5);
  assign w695[41] = |(datain[147:144] ^ 9);
  assign w695[42] = |(datain[143:140] ^ 0);
  assign w695[43] = |(datain[139:136] ^ 3);
  assign w695[44] = |(datain[135:132] ^ 12);
  assign w695[45] = |(datain[131:128] ^ 10);
  assign w695[46] = |(datain[127:124] ^ 5);
  assign w695[47] = |(datain[123:120] ^ 10);
  assign w695[48] = |(datain[119:116] ^ 11);
  assign w695[49] = |(datain[115:112] ^ 4);
  assign w695[50] = |(datain[111:108] ^ 4);
  assign w695[51] = |(datain[107:104] ^ 0);
  assign w695[52] = |(datain[103:100] ^ 12);
  assign w695[53] = |(datain[99:96] ^ 13);
  assign w695[54] = |(datain[95:92] ^ 2);
  assign w695[55] = |(datain[91:88] ^ 1);
  assign w695[56] = |(datain[87:84] ^ 7);
  assign w695[57] = |(datain[83:80] ^ 2);
  assign w695[58] = |(datain[79:76] ^ 1);
  assign w695[59] = |(datain[75:72] ^ 3);
  assign w695[60] = |(datain[71:68] ^ 11);
  assign w695[61] = |(datain[67:64] ^ 8);
  assign w695[62] = |(datain[63:60] ^ 0);
  assign w695[63] = |(datain[59:56] ^ 0);
  assign w695[64] = |(datain[55:52] ^ 4);
  assign w695[65] = |(datain[51:48] ^ 2);
  assign w695[66] = |(datain[47:44] ^ 9);
  assign w695[67] = |(datain[43:40] ^ 9);
  assign w695[68] = |(datain[39:36] ^ 3);
  assign w695[69] = |(datain[35:32] ^ 3);
  assign w695[70] = |(datain[31:28] ^ 12);
  assign w695[71] = |(datain[27:24] ^ 9);
  assign w695[72] = |(datain[23:20] ^ 12);
  assign w695[73] = |(datain[19:16] ^ 13);
  assign w695[74] = |(datain[15:12] ^ 2);
  assign w695[75] = |(datain[11:8] ^ 1);
  assign comp[695] = ~(|w695);
  wire [76-1:0] w696;
  assign w696[0] = |(datain[311:308] ^ 12);
  assign w696[1] = |(datain[307:304] ^ 13);
  assign w696[2] = |(datain[303:300] ^ 2);
  assign w696[3] = |(datain[299:296] ^ 1);
  assign w696[4] = |(datain[295:292] ^ 2);
  assign w696[5] = |(datain[291:288] ^ 14);
  assign w696[6] = |(datain[287:284] ^ 10);
  assign w696[7] = |(datain[283:280] ^ 3);
  assign w696[8] = |(datain[279:276] ^ 11);
  assign w696[9] = |(datain[275:272] ^ 9);
  assign w696[10] = |(datain[271:268] ^ 0);
  assign w696[11] = |(datain[267:264] ^ 1);
  assign w696[12] = |(datain[263:260] ^ 11);
  assign w696[13] = |(datain[259:256] ^ 4);
  assign w696[14] = |(datain[255:252] ^ 4);
  assign w696[15] = |(datain[251:248] ^ 0);
  assign w696[16] = |(datain[247:244] ^ 11);
  assign w696[17] = |(datain[243:240] ^ 9);
  assign w696[18] = |(datain[239:236] ^ 13);
  assign w696[19] = |(datain[235:232] ^ 13);
  assign w696[20] = |(datain[231:228] ^ 0);
  assign w696[21] = |(datain[227:224] ^ 1);
  assign w696[22] = |(datain[223:220] ^ 3);
  assign w696[23] = |(datain[219:216] ^ 3);
  assign w696[24] = |(datain[215:212] ^ 13);
  assign w696[25] = |(datain[211:208] ^ 2);
  assign w696[26] = |(datain[207:204] ^ 12);
  assign w696[27] = |(datain[203:200] ^ 13);
  assign w696[28] = |(datain[199:196] ^ 2);
  assign w696[29] = |(datain[195:192] ^ 1);
  assign w696[30] = |(datain[191:188] ^ 3);
  assign w696[31] = |(datain[187:184] ^ 3);
  assign w696[32] = |(datain[183:180] ^ 12);
  assign w696[33] = |(datain[179:176] ^ 9);
  assign w696[34] = |(datain[175:172] ^ 3);
  assign w696[35] = |(datain[171:168] ^ 3);
  assign w696[36] = |(datain[167:164] ^ 13);
  assign w696[37] = |(datain[163:160] ^ 2);
  assign w696[38] = |(datain[159:156] ^ 11);
  assign w696[39] = |(datain[155:152] ^ 8);
  assign w696[40] = |(datain[151:148] ^ 0);
  assign w696[41] = |(datain[147:144] ^ 0);
  assign w696[42] = |(datain[143:140] ^ 4);
  assign w696[43] = |(datain[139:136] ^ 2);
  assign w696[44] = |(datain[135:132] ^ 12);
  assign w696[45] = |(datain[131:128] ^ 13);
  assign w696[46] = |(datain[127:124] ^ 2);
  assign w696[47] = |(datain[123:120] ^ 1);
  assign w696[48] = |(datain[119:116] ^ 11);
  assign w696[49] = |(datain[115:112] ^ 4);
  assign w696[50] = |(datain[111:108] ^ 4);
  assign w696[51] = |(datain[107:104] ^ 0);
  assign w696[52] = |(datain[103:100] ^ 11);
  assign w696[53] = |(datain[99:96] ^ 9);
  assign w696[54] = |(datain[95:92] ^ 0);
  assign w696[55] = |(datain[91:88] ^ 3);
  assign w696[56] = |(datain[87:84] ^ 0);
  assign w696[57] = |(datain[83:80] ^ 0);
  assign w696[58] = |(datain[79:76] ^ 11);
  assign w696[59] = |(datain[75:72] ^ 10);
  assign w696[60] = |(datain[71:68] ^ 11);
  assign w696[61] = |(datain[67:64] ^ 8);
  assign w696[62] = |(datain[63:60] ^ 0);
  assign w696[63] = |(datain[59:56] ^ 1);
  assign w696[64] = |(datain[55:52] ^ 12);
  assign w696[65] = |(datain[51:48] ^ 13);
  assign w696[66] = |(datain[47:44] ^ 2);
  assign w696[67] = |(datain[43:40] ^ 1);
  assign w696[68] = |(datain[39:36] ^ 11);
  assign w696[69] = |(datain[35:32] ^ 8);
  assign w696[70] = |(datain[31:28] ^ 0);
  assign w696[71] = |(datain[27:24] ^ 1);
  assign w696[72] = |(datain[23:20] ^ 5);
  assign w696[73] = |(datain[19:16] ^ 7);
  assign w696[74] = |(datain[15:12] ^ 2);
  assign w696[75] = |(datain[11:8] ^ 14);
  assign comp[696] = ~(|w696);
  wire [46-1:0] w697;
  assign w697[0] = |(datain[311:308] ^ 11);
  assign w697[1] = |(datain[307:304] ^ 9);
  assign w697[2] = |(datain[303:300] ^ 2);
  assign w697[3] = |(datain[299:296] ^ 3);
  assign w697[4] = |(datain[295:292] ^ 0);
  assign w697[5] = |(datain[291:288] ^ 9);
  assign w697[6] = |(datain[287:284] ^ 0);
  assign w697[7] = |(datain[283:280] ^ 15);
  assign w697[8] = |(datain[279:276] ^ 4);
  assign w697[9] = |(datain[275:272] ^ 11);
  assign w697[10] = |(datain[271:268] ^ 8);
  assign w697[11] = |(datain[267:264] ^ 14);
  assign w697[12] = |(datain[263:260] ^ 6);
  assign w697[13] = |(datain[259:256] ^ 14);
  assign w697[14] = |(datain[255:252] ^ 7);
  assign w697[15] = |(datain[251:248] ^ 11);
  assign w697[16] = |(datain[247:244] ^ 3);
  assign w697[17] = |(datain[243:240] ^ 5);
  assign w697[18] = |(datain[239:236] ^ 8);
  assign w697[19] = |(datain[235:232] ^ 12);
  assign w697[20] = |(datain[231:228] ^ 8);
  assign w697[21] = |(datain[227:224] ^ 13);
  assign w697[22] = |(datain[223:220] ^ 3);
  assign w697[23] = |(datain[219:216] ^ 3);
  assign w697[24] = |(datain[215:212] ^ 9);
  assign w697[25] = |(datain[211:208] ^ 12);
  assign w697[26] = |(datain[207:204] ^ 10);
  assign w697[27] = |(datain[203:200] ^ 4);
  assign w697[28] = |(datain[199:196] ^ 0);
  assign w697[29] = |(datain[195:192] ^ 13);
  assign w697[30] = |(datain[191:188] ^ 11);
  assign w697[31] = |(datain[187:184] ^ 9);
  assign w697[32] = |(datain[183:180] ^ 3);
  assign w697[33] = |(datain[179:176] ^ 14);
  assign w697[34] = |(datain[175:172] ^ 7);
  assign w697[35] = |(datain[171:168] ^ 0);
  assign w697[36] = |(datain[167:164] ^ 0);
  assign w697[37] = |(datain[163:160] ^ 15);
  assign w697[38] = |(datain[159:156] ^ 4);
  assign w697[39] = |(datain[155:152] ^ 11);
  assign w697[40] = |(datain[151:148] ^ 8);
  assign w697[41] = |(datain[147:144] ^ 14);
  assign w697[42] = |(datain[143:140] ^ 6);
  assign w697[43] = |(datain[139:136] ^ 14);
  assign w697[44] = |(datain[135:132] ^ 7);
  assign w697[45] = |(datain[131:128] ^ 11);
  assign comp[697] = ~(|w697);
  wire [76-1:0] w698;
  assign w698[0] = |(datain[311:308] ^ 2);
  assign w698[1] = |(datain[307:304] ^ 4);
  assign w698[2] = |(datain[303:300] ^ 8);
  assign w698[3] = |(datain[299:296] ^ 3);
  assign w698[4] = |(datain[295:292] ^ 3);
  assign w698[5] = |(datain[291:288] ^ 14);
  assign w698[6] = |(datain[287:284] ^ 9);
  assign w698[7] = |(datain[283:280] ^ 12);
  assign w698[8] = |(datain[279:276] ^ 0);
  assign w698[9] = |(datain[275:272] ^ 0);
  assign w698[10] = |(datain[271:268] ^ 0);
  assign w698[11] = |(datain[267:264] ^ 0);
  assign w698[12] = |(datain[263:260] ^ 7);
  assign w698[13] = |(datain[259:256] ^ 5);
  assign w698[14] = |(datain[255:252] ^ 1);
  assign w698[15] = |(datain[251:248] ^ 7);
  assign w698[16] = |(datain[247:244] ^ 11);
  assign w698[17] = |(datain[243:240] ^ 10);
  assign w698[18] = |(datain[239:236] ^ 9);
  assign w698[19] = |(datain[235:232] ^ 14);
  assign w698[20] = |(datain[231:228] ^ 0);
  assign w698[21] = |(datain[227:224] ^ 0);
  assign w698[22] = |(datain[223:220] ^ 11);
  assign w698[23] = |(datain[219:216] ^ 8);
  assign w698[24] = |(datain[215:212] ^ 0);
  assign w698[25] = |(datain[211:208] ^ 1);
  assign w698[26] = |(datain[207:204] ^ 3);
  assign w698[27] = |(datain[203:200] ^ 13);
  assign w698[28] = |(datain[199:196] ^ 12);
  assign w698[29] = |(datain[195:192] ^ 13);
  assign w698[30] = |(datain[191:188] ^ 2);
  assign w698[31] = |(datain[187:184] ^ 1);
  assign w698[32] = |(datain[183:180] ^ 9);
  assign w698[33] = |(datain[179:176] ^ 3);
  assign w698[34] = |(datain[175:172] ^ 11);
  assign w698[35] = |(datain[171:168] ^ 4);
  assign w698[36] = |(datain[167:164] ^ 4);
  assign w698[37] = |(datain[163:160] ^ 0);
  assign w698[38] = |(datain[159:156] ^ 11);
  assign w698[39] = |(datain[155:152] ^ 10);
  assign w698[40] = |(datain[151:148] ^ 0);
  assign w698[41] = |(datain[147:144] ^ 0);
  assign w698[42] = |(datain[143:140] ^ 0);
  assign w698[43] = |(datain[139:136] ^ 1);
  assign w698[44] = |(datain[135:132] ^ 11);
  assign w698[45] = |(datain[131:128] ^ 9);
  assign w698[46] = |(datain[127:124] ^ 9);
  assign w698[47] = |(datain[123:120] ^ 12);
  assign w698[48] = |(datain[119:116] ^ 0);
  assign w698[49] = |(datain[115:112] ^ 0);
  assign w698[50] = |(datain[111:108] ^ 12);
  assign w698[51] = |(datain[107:104] ^ 13);
  assign w698[52] = |(datain[103:100] ^ 2);
  assign w698[53] = |(datain[99:96] ^ 1);
  assign w698[54] = |(datain[95:92] ^ 11);
  assign w698[55] = |(datain[91:88] ^ 4);
  assign w698[56] = |(datain[87:84] ^ 3);
  assign w698[57] = |(datain[83:80] ^ 14);
  assign w698[58] = |(datain[79:76] ^ 12);
  assign w698[59] = |(datain[75:72] ^ 13);
  assign w698[60] = |(datain[71:68] ^ 2);
  assign w698[61] = |(datain[67:64] ^ 1);
  assign w698[62] = |(datain[63:60] ^ 11);
  assign w698[63] = |(datain[59:56] ^ 4);
  assign w698[64] = |(datain[55:52] ^ 4);
  assign w698[65] = |(datain[51:48] ^ 15);
  assign w698[66] = |(datain[47:44] ^ 12);
  assign w698[67] = |(datain[43:40] ^ 13);
  assign w698[68] = |(datain[39:36] ^ 2);
  assign w698[69] = |(datain[35:32] ^ 1);
  assign w698[70] = |(datain[31:28] ^ 7);
  assign w698[71] = |(datain[27:24] ^ 3);
  assign w698[72] = |(datain[23:20] ^ 13);
  assign w698[73] = |(datain[19:16] ^ 10);
  assign w698[74] = |(datain[15:12] ^ 12);
  assign w698[75] = |(datain[11:8] ^ 3);
  assign comp[698] = ~(|w698);
  wire [74-1:0] w699;
  assign w699[0] = |(datain[311:308] ^ 3);
  assign w699[1] = |(datain[307:304] ^ 3);
  assign w699[2] = |(datain[303:300] ^ 12);
  assign w699[3] = |(datain[299:296] ^ 9);
  assign w699[4] = |(datain[295:292] ^ 9);
  assign w699[5] = |(datain[291:288] ^ 9);
  assign w699[6] = |(datain[287:284] ^ 12);
  assign w699[7] = |(datain[283:280] ^ 13);
  assign w699[8] = |(datain[279:276] ^ 2);
  assign w699[9] = |(datain[275:272] ^ 1);
  assign w699[10] = |(datain[271:268] ^ 11);
  assign w699[11] = |(datain[267:264] ^ 4);
  assign w699[12] = |(datain[263:260] ^ 4);
  assign w699[13] = |(datain[259:256] ^ 0);
  assign w699[14] = |(datain[255:252] ^ 8);
  assign w699[15] = |(datain[251:248] ^ 11);
  assign w699[16] = |(datain[247:244] ^ 13);
  assign w699[17] = |(datain[243:240] ^ 6);
  assign w699[18] = |(datain[239:236] ^ 11);
  assign w699[19] = |(datain[235:232] ^ 9);
  assign w699[20] = |(datain[231:228] ^ 1);
  assign w699[21] = |(datain[227:224] ^ 12);
  assign w699[22] = |(datain[223:220] ^ 0);
  assign w699[23] = |(datain[219:216] ^ 0);
  assign w699[24] = |(datain[215:212] ^ 12);
  assign w699[25] = |(datain[211:208] ^ 13);
  assign w699[26] = |(datain[207:204] ^ 2);
  assign w699[27] = |(datain[203:200] ^ 1);
  assign w699[28] = |(datain[199:196] ^ 11);
  assign w699[29] = |(datain[195:192] ^ 8);
  assign w699[30] = |(datain[191:188] ^ 0);
  assign w699[31] = |(datain[187:184] ^ 2);
  assign w699[32] = |(datain[183:180] ^ 4);
  assign w699[33] = |(datain[179:176] ^ 2);
  assign w699[34] = |(datain[175:172] ^ 9);
  assign w699[35] = |(datain[171:168] ^ 9);
  assign w699[36] = |(datain[167:164] ^ 3);
  assign w699[37] = |(datain[163:160] ^ 3);
  assign w699[38] = |(datain[159:156] ^ 12);
  assign w699[39] = |(datain[155:152] ^ 9);
  assign w699[40] = |(datain[151:148] ^ 12);
  assign w699[41] = |(datain[147:144] ^ 13);
  assign w699[42] = |(datain[143:140] ^ 2);
  assign w699[43] = |(datain[139:136] ^ 1);
  assign w699[44] = |(datain[135:132] ^ 1);
  assign w699[45] = |(datain[131:128] ^ 14);
  assign w699[46] = |(datain[127:124] ^ 0);
  assign w699[47] = |(datain[123:120] ^ 7);
  assign w699[48] = |(datain[119:116] ^ 11);
  assign w699[49] = |(datain[115:112] ^ 14);
  assign w699[50] = |(datain[111:108] ^ 8);
  assign w699[51] = |(datain[107:104] ^ 4);
  assign w699[52] = |(datain[103:100] ^ 0);
  assign w699[53] = |(datain[99:96] ^ 3);
  assign w699[54] = |(datain[95:92] ^ 11);
  assign w699[55] = |(datain[91:88] ^ 15);
  assign w699[56] = |(datain[87:84] ^ 0);
  assign w699[57] = |(datain[83:80] ^ 5);
  assign w699[58] = |(datain[79:76] ^ 0);
  assign w699[59] = |(datain[75:72] ^ 0);
  assign w699[60] = |(datain[71:68] ^ 14);
  assign w699[61] = |(datain[67:64] ^ 4);
  assign w699[62] = |(datain[63:60] ^ 4);
  assign w699[63] = |(datain[59:56] ^ 0);
  assign w699[64] = |(datain[55:52] ^ 11);
  assign w699[65] = |(datain[51:48] ^ 10);
  assign w699[66] = |(datain[47:44] ^ 0);
  assign w699[67] = |(datain[43:40] ^ 3);
  assign w699[68] = |(datain[39:36] ^ 0);
  assign w699[69] = |(datain[35:32] ^ 0);
  assign w699[70] = |(datain[31:28] ^ 2);
  assign w699[71] = |(datain[27:24] ^ 3);
  assign w699[72] = |(datain[23:20] ^ 12);
  assign w699[73] = |(datain[19:16] ^ 2);
  assign comp[699] = ~(|w699);
  wire [36-1:0] w700;
  assign w700[0] = |(datain[311:308] ^ 11);
  assign w700[1] = |(datain[307:304] ^ 8);
  assign w700[2] = |(datain[303:300] ^ 12);
  assign w700[3] = |(datain[299:296] ^ 10);
  assign w700[4] = |(datain[295:292] ^ 0);
  assign w700[5] = |(datain[291:288] ^ 0);
  assign w700[6] = |(datain[287:284] ^ 5);
  assign w700[7] = |(datain[283:280] ^ 0);
  assign w700[8] = |(datain[279:276] ^ 12);
  assign w700[9] = |(datain[275:272] ^ 11);
  assign w700[10] = |(datain[271:268] ^ 3);
  assign w700[11] = |(datain[267:264] ^ 1);
  assign w700[12] = |(datain[263:260] ^ 12);
  assign w700[13] = |(datain[259:256] ^ 0);
  assign w700[14] = |(datain[255:252] ^ 12);
  assign w700[15] = |(datain[251:248] ^ 13);
  assign w700[16] = |(datain[247:244] ^ 1);
  assign w700[17] = |(datain[243:240] ^ 3);
  assign w700[18] = |(datain[239:236] ^ 3);
  assign w700[19] = |(datain[235:232] ^ 1);
  assign w700[20] = |(datain[231:228] ^ 12);
  assign w700[21] = |(datain[227:224] ^ 0);
  assign w700[22] = |(datain[223:220] ^ 8);
  assign w700[23] = |(datain[219:216] ^ 14);
  assign w700[24] = |(datain[215:212] ^ 12);
  assign w700[25] = |(datain[211:208] ^ 0);
  assign w700[26] = |(datain[207:204] ^ 11);
  assign w700[27] = |(datain[203:200] ^ 8);
  assign w700[28] = |(datain[199:196] ^ 0);
  assign w700[29] = |(datain[195:192] ^ 1);
  assign w700[30] = |(datain[191:188] ^ 0);
  assign w700[31] = |(datain[187:184] ^ 2);
  assign w700[32] = |(datain[183:180] ^ 11);
  assign w700[33] = |(datain[179:176] ^ 11);
  assign w700[34] = |(datain[175:172] ^ 0);
  assign w700[35] = |(datain[171:168] ^ 0);
  assign comp[700] = ~(|w700);
  wire [32-1:0] w701;
  assign w701[0] = |(datain[311:308] ^ 11);
  assign w701[1] = |(datain[307:304] ^ 9);
  assign w701[2] = |(datain[303:300] ^ 0);
  assign w701[3] = |(datain[299:296] ^ 8);
  assign w701[4] = |(datain[295:292] ^ 2);
  assign w701[5] = |(datain[291:288] ^ 7);
  assign w701[6] = |(datain[287:284] ^ 11);
  assign w701[7] = |(datain[283:280] ^ 10);
  assign w701[8] = |(datain[279:276] ^ 0);
  assign w701[9] = |(datain[275:272] ^ 0);
  assign w701[10] = |(datain[271:268] ^ 0);
  assign w701[11] = |(datain[267:264] ^ 1);
  assign w701[12] = |(datain[263:260] ^ 12);
  assign w701[13] = |(datain[259:256] ^ 13);
  assign w701[14] = |(datain[255:252] ^ 1);
  assign w701[15] = |(datain[251:248] ^ 3);
  assign w701[16] = |(datain[247:244] ^ 7);
  assign w701[17] = |(datain[243:240] ^ 2);
  assign w701[18] = |(datain[239:236] ^ 15);
  assign w701[19] = |(datain[235:232] ^ 1);
  assign w701[20] = |(datain[231:228] ^ 0);
  assign w701[21] = |(datain[227:224] ^ 14);
  assign w701[22] = |(datain[223:220] ^ 0);
  assign w701[23] = |(datain[219:216] ^ 7);
  assign w701[24] = |(datain[215:212] ^ 11);
  assign w701[25] = |(datain[211:208] ^ 8);
  assign w701[26] = |(datain[207:204] ^ 0);
  assign w701[27] = |(datain[203:200] ^ 1);
  assign w701[28] = |(datain[199:196] ^ 0);
  assign w701[29] = |(datain[195:192] ^ 2);
  assign w701[30] = |(datain[191:188] ^ 11);
  assign w701[31] = |(datain[187:184] ^ 11);
  assign comp[701] = ~(|w701);
  wire [42-1:0] w702;
  assign w702[0] = |(datain[311:308] ^ 4);
  assign w702[1] = |(datain[307:304] ^ 2);
  assign w702[2] = |(datain[303:300] ^ 4);
  assign w702[3] = |(datain[299:296] ^ 1);
  assign w702[4] = |(datain[295:292] ^ 7);
  assign w702[5] = |(datain[291:288] ^ 4);
  assign w702[6] = |(datain[287:284] ^ 4);
  assign w702[7] = |(datain[283:280] ^ 1);
  assign w702[8] = |(datain[279:276] ^ 11);
  assign w702[9] = |(datain[275:272] ^ 11);
  assign w702[10] = |(datain[271:268] ^ 8);
  assign w702[11] = |(datain[267:264] ^ 0);
  assign w702[12] = |(datain[263:260] ^ 0);
  assign w702[13] = |(datain[259:256] ^ 0);
  assign w702[14] = |(datain[255:252] ^ 8);
  assign w702[15] = |(datain[251:248] ^ 11);
  assign w702[16] = |(datain[247:244] ^ 5);
  assign w702[17] = |(datain[243:240] ^ 7);
  assign w702[18] = |(datain[239:236] ^ 1);
  assign w702[19] = |(datain[235:232] ^ 10);
  assign w702[20] = |(datain[231:228] ^ 8);
  assign w702[21] = |(datain[227:224] ^ 1);
  assign w702[22] = |(datain[223:220] ^ 12);
  assign w702[23] = |(datain[219:216] ^ 2);
  assign w702[24] = |(datain[215:212] ^ 11);
  assign w702[25] = |(datain[211:208] ^ 5);
  assign w702[26] = |(datain[207:204] ^ 0);
  assign w702[27] = |(datain[203:200] ^ 0);
  assign w702[28] = |(datain[199:196] ^ 8);
  assign w702[29] = |(datain[195:192] ^ 1);
  assign w702[30] = |(datain[191:188] ^ 12);
  assign w702[31] = |(datain[187:184] ^ 2);
  assign w702[32] = |(datain[183:180] ^ 0);
  assign w702[33] = |(datain[179:176] ^ 0);
  assign w702[34] = |(datain[175:172] ^ 0);
  assign w702[35] = |(datain[171:168] ^ 1);
  assign w702[36] = |(datain[167:164] ^ 8);
  assign w702[37] = |(datain[163:160] ^ 9);
  assign w702[38] = |(datain[159:156] ^ 1);
  assign w702[39] = |(datain[155:152] ^ 6);
  assign w702[40] = |(datain[151:148] ^ 0);
  assign w702[41] = |(datain[147:144] ^ 6);
  assign comp[702] = ~(|w702);
  wire [44-1:0] w703;
  assign w703[0] = |(datain[311:308] ^ 0);
  assign w703[1] = |(datain[307:304] ^ 1);
  assign w703[2] = |(datain[303:300] ^ 8);
  assign w703[3] = |(datain[299:296] ^ 1);
  assign w703[4] = |(datain[295:292] ^ 12);
  assign w703[5] = |(datain[291:288] ^ 6);
  assign w703[6] = |(datain[287:284] ^ 4);
  assign w703[7] = |(datain[283:280] ^ 6);
  assign w703[8] = |(datain[279:276] ^ 0);
  assign w703[9] = |(datain[275:272] ^ 1);
  assign w703[10] = |(datain[271:268] ^ 11);
  assign w703[11] = |(datain[267:264] ^ 9);
  assign w703[12] = |(datain[263:260] ^ 0);
  assign w703[13] = |(datain[259:256] ^ 4);
  assign w703[14] = |(datain[255:252] ^ 0);
  assign w703[15] = |(datain[251:248] ^ 0);
  assign w703[16] = |(datain[247:244] ^ 15);
  assign w703[17] = |(datain[243:240] ^ 12);
  assign w703[18] = |(datain[239:236] ^ 15);
  assign w703[19] = |(datain[235:232] ^ 3);
  assign w703[20] = |(datain[231:228] ^ 10);
  assign w703[21] = |(datain[227:224] ^ 4);
  assign w703[22] = |(datain[223:220] ^ 5);
  assign w703[23] = |(datain[219:216] ^ 14);
  assign w703[24] = |(datain[215:212] ^ 11);
  assign w703[25] = |(datain[211:208] ^ 8);
  assign w703[26] = |(datain[207:204] ^ 11);
  assign w703[27] = |(datain[203:200] ^ 10);
  assign w703[28] = |(datain[199:196] ^ 11);
  assign w703[29] = |(datain[195:192] ^ 10);
  assign w703[30] = |(datain[191:188] ^ 12);
  assign w703[31] = |(datain[187:184] ^ 13);
  assign w703[32] = |(datain[183:180] ^ 2);
  assign w703[33] = |(datain[179:176] ^ 1);
  assign w703[34] = |(datain[175:172] ^ 3);
  assign w703[35] = |(datain[171:168] ^ 13);
  assign w703[36] = |(datain[167:164] ^ 12);
  assign w703[37] = |(datain[163:160] ^ 12);
  assign w703[38] = |(datain[159:156] ^ 15);
  assign w703[39] = |(datain[155:152] ^ 10);
  assign w703[40] = |(datain[151:148] ^ 7);
  assign w703[41] = |(datain[147:144] ^ 5);
  assign w703[42] = |(datain[143:140] ^ 0);
  assign w703[43] = |(datain[139:136] ^ 3);
  assign comp[703] = ~(|w703);
  wire [76-1:0] w704;
  assign w704[0] = |(datain[311:308] ^ 8);
  assign w704[1] = |(datain[307:304] ^ 12);
  assign w704[2] = |(datain[303:300] ^ 12);
  assign w704[3] = |(datain[299:296] ^ 8);
  assign w704[4] = |(datain[295:292] ^ 8);
  assign w704[5] = |(datain[291:288] ^ 14);
  assign w704[6] = |(datain[287:284] ^ 13);
  assign w704[7] = |(datain[283:280] ^ 8);
  assign w704[8] = |(datain[279:276] ^ 11);
  assign w704[9] = |(datain[275:272] ^ 4);
  assign w704[10] = |(datain[271:268] ^ 4);
  assign w704[11] = |(datain[267:264] ^ 0);
  assign w704[12] = |(datain[263:260] ^ 3);
  assign w704[13] = |(datain[259:256] ^ 3);
  assign w704[14] = |(datain[255:252] ^ 13);
  assign w704[15] = |(datain[251:248] ^ 2);
  assign w704[16] = |(datain[247:244] ^ 11);
  assign w704[17] = |(datain[243:240] ^ 9);
  assign w704[18] = |(datain[239:236] ^ 6);
  assign w704[19] = |(datain[235:232] ^ 4);
  assign w704[20] = |(datain[231:228] ^ 0);
  assign w704[21] = |(datain[227:224] ^ 1);
  assign w704[22] = |(datain[223:220] ^ 9);
  assign w704[23] = |(datain[219:216] ^ 0);
  assign w704[24] = |(datain[215:212] ^ 12);
  assign w704[25] = |(datain[211:208] ^ 13);
  assign w704[26] = |(datain[207:204] ^ 2);
  assign w704[27] = |(datain[203:200] ^ 1);
  assign w704[28] = |(datain[199:196] ^ 3);
  assign w704[29] = |(datain[195:192] ^ 3);
  assign w704[30] = |(datain[191:188] ^ 12);
  assign w704[31] = |(datain[187:184] ^ 9);
  assign w704[32] = |(datain[183:180] ^ 3);
  assign w704[33] = |(datain[179:176] ^ 3);
  assign w704[34] = |(datain[175:172] ^ 13);
  assign w704[35] = |(datain[171:168] ^ 2);
  assign w704[36] = |(datain[167:164] ^ 11);
  assign w704[37] = |(datain[163:160] ^ 8);
  assign w704[38] = |(datain[159:156] ^ 0);
  assign w704[39] = |(datain[155:152] ^ 0);
  assign w704[40] = |(datain[151:148] ^ 4);
  assign w704[41] = |(datain[147:144] ^ 2);
  assign w704[42] = |(datain[143:140] ^ 12);
  assign w704[43] = |(datain[139:136] ^ 13);
  assign w704[44] = |(datain[135:132] ^ 2);
  assign w704[45] = |(datain[131:128] ^ 1);
  assign w704[46] = |(datain[127:124] ^ 11);
  assign w704[47] = |(datain[123:120] ^ 4);
  assign w704[48] = |(datain[119:116] ^ 4);
  assign w704[49] = |(datain[115:112] ^ 0);
  assign w704[50] = |(datain[111:108] ^ 11);
  assign w704[51] = |(datain[107:104] ^ 10);
  assign w704[52] = |(datain[103:100] ^ 5);
  assign w704[53] = |(datain[99:96] ^ 1);
  assign w704[54] = |(datain[95:92] ^ 0);
  assign w704[55] = |(datain[91:88] ^ 1);
  assign w704[56] = |(datain[87:84] ^ 11);
  assign w704[57] = |(datain[83:80] ^ 9);
  assign w704[58] = |(datain[79:76] ^ 0);
  assign w704[59] = |(datain[75:72] ^ 4);
  assign w704[60] = |(datain[71:68] ^ 0);
  assign w704[61] = |(datain[67:64] ^ 0);
  assign w704[62] = |(datain[63:60] ^ 12);
  assign w704[63] = |(datain[59:56] ^ 13);
  assign w704[64] = |(datain[55:52] ^ 2);
  assign w704[65] = |(datain[51:48] ^ 1);
  assign w704[66] = |(datain[47:44] ^ 11);
  assign w704[67] = |(datain[43:40] ^ 4);
  assign w704[68] = |(datain[39:36] ^ 3);
  assign w704[69] = |(datain[35:32] ^ 14);
  assign w704[70] = |(datain[31:28] ^ 12);
  assign w704[71] = |(datain[27:24] ^ 13);
  assign w704[72] = |(datain[23:20] ^ 2);
  assign w704[73] = |(datain[19:16] ^ 1);
  assign w704[74] = |(datain[15:12] ^ 5);
  assign w704[75] = |(datain[11:8] ^ 10);
  assign comp[704] = ~(|w704);
  wire [74-1:0] w705;
  assign w705[0] = |(datain[311:308] ^ 7);
  assign w705[1] = |(datain[307:304] ^ 12);
  assign w705[2] = |(datain[303:300] ^ 6);
  assign w705[3] = |(datain[299:296] ^ 3);
  assign w705[4] = |(datain[295:292] ^ 3);
  assign w705[5] = |(datain[291:288] ^ 13);
  assign w705[6] = |(datain[287:284] ^ 0);
  assign w705[7] = |(datain[283:280] ^ 0);
  assign w705[8] = |(datain[279:276] ^ 15);
  assign w705[9] = |(datain[275:272] ^ 10);
  assign w705[10] = |(datain[271:268] ^ 7);
  assign w705[11] = |(datain[267:264] ^ 7);
  assign w705[12] = |(datain[263:260] ^ 5);
  assign w705[13] = |(datain[259:256] ^ 14);
  assign w705[14] = |(datain[255:252] ^ 2);
  assign w705[15] = |(datain[251:248] ^ 13);
  assign w705[16] = |(datain[247:244] ^ 0);
  assign w705[17] = |(datain[243:240] ^ 3);
  assign w705[18] = |(datain[239:236] ^ 0);
  assign w705[19] = |(datain[235:232] ^ 0);
  assign w705[20] = |(datain[231:228] ^ 2);
  assign w705[21] = |(datain[227:224] ^ 14);
  assign w705[22] = |(datain[223:220] ^ 10);
  assign w705[23] = |(datain[219:216] ^ 3);
  assign w705[24] = |(datain[215:212] ^ 9);
  assign w705[25] = |(datain[211:208] ^ 10);
  assign w705[26] = |(datain[207:204] ^ 0);
  assign w705[27] = |(datain[203:200] ^ 1);
  assign w705[28] = |(datain[199:196] ^ 2);
  assign w705[29] = |(datain[195:192] ^ 14);
  assign w705[30] = |(datain[191:188] ^ 8);
  assign w705[31] = |(datain[187:184] ^ 0);
  assign w705[32] = |(datain[183:180] ^ 3);
  assign w705[33] = |(datain[179:176] ^ 14);
  assign w705[34] = |(datain[175:172] ^ 9);
  assign w705[35] = |(datain[171:168] ^ 8);
  assign w705[36] = |(datain[167:164] ^ 0);
  assign w705[37] = |(datain[163:160] ^ 1);
  assign w705[38] = |(datain[159:156] ^ 0);
  assign w705[39] = |(datain[155:152] ^ 15);
  assign w705[40] = |(datain[151:148] ^ 7);
  assign w705[41] = |(datain[147:144] ^ 4);
  assign w705[42] = |(datain[143:140] ^ 4);
  assign w705[43] = |(datain[139:136] ^ 15);
  assign w705[44] = |(datain[135:132] ^ 8);
  assign w705[45] = |(datain[131:128] ^ 12);
  assign w705[46] = |(datain[127:124] ^ 12);
  assign w705[47] = |(datain[123:120] ^ 8);
  assign w705[48] = |(datain[119:116] ^ 8);
  assign w705[49] = |(datain[115:112] ^ 14);
  assign w705[50] = |(datain[111:108] ^ 13);
  assign w705[51] = |(datain[107:104] ^ 8);
  assign w705[52] = |(datain[103:100] ^ 11);
  assign w705[53] = |(datain[99:96] ^ 4);
  assign w705[54] = |(datain[95:92] ^ 4);
  assign w705[55] = |(datain[91:88] ^ 0);
  assign w705[56] = |(datain[87:84] ^ 3);
  assign w705[57] = |(datain[83:80] ^ 3);
  assign w705[58] = |(datain[79:76] ^ 13);
  assign w705[59] = |(datain[75:72] ^ 2);
  assign w705[60] = |(datain[71:68] ^ 11);
  assign w705[61] = |(datain[67:64] ^ 9);
  assign w705[62] = |(datain[63:60] ^ 10);
  assign w705[63] = |(datain[59:56] ^ 13);
  assign w705[64] = |(datain[55:52] ^ 0);
  assign w705[65] = |(datain[51:48] ^ 1);
  assign w705[66] = |(datain[47:44] ^ 12);
  assign w705[67] = |(datain[43:40] ^ 13);
  assign w705[68] = |(datain[39:36] ^ 2);
  assign w705[69] = |(datain[35:32] ^ 1);
  assign w705[70] = |(datain[31:28] ^ 3);
  assign w705[71] = |(datain[27:24] ^ 3);
  assign w705[72] = |(datain[23:20] ^ 12);
  assign w705[73] = |(datain[19:16] ^ 9);
  assign comp[705] = ~(|w705);
  wire [46-1:0] w706;
  assign w706[0] = |(datain[311:308] ^ 13);
  assign w706[1] = |(datain[307:304] ^ 8);
  assign w706[2] = |(datain[303:300] ^ 11);
  assign w706[3] = |(datain[299:296] ^ 4);
  assign w706[4] = |(datain[295:292] ^ 4);
  assign w706[5] = |(datain[291:288] ^ 0);
  assign w706[6] = |(datain[287:284] ^ 3);
  assign w706[7] = |(datain[283:280] ^ 3);
  assign w706[8] = |(datain[279:276] ^ 13);
  assign w706[9] = |(datain[275:272] ^ 2);
  assign w706[10] = |(datain[271:268] ^ 11);
  assign w706[11] = |(datain[267:264] ^ 9);
  assign w706[12] = |(datain[263:260] ^ 13);
  assign w706[13] = |(datain[259:256] ^ 6);
  assign w706[14] = |(datain[255:252] ^ 0);
  assign w706[15] = |(datain[251:248] ^ 1);
  assign w706[16] = |(datain[247:244] ^ 12);
  assign w706[17] = |(datain[243:240] ^ 13);
  assign w706[18] = |(datain[239:236] ^ 2);
  assign w706[19] = |(datain[235:232] ^ 1);
  assign w706[20] = |(datain[231:228] ^ 3);
  assign w706[21] = |(datain[227:224] ^ 3);
  assign w706[22] = |(datain[223:220] ^ 12);
  assign w706[23] = |(datain[219:216] ^ 9);
  assign w706[24] = |(datain[215:212] ^ 3);
  assign w706[25] = |(datain[211:208] ^ 3);
  assign w706[26] = |(datain[207:204] ^ 13);
  assign w706[27] = |(datain[203:200] ^ 2);
  assign w706[28] = |(datain[199:196] ^ 11);
  assign w706[29] = |(datain[195:192] ^ 8);
  assign w706[30] = |(datain[191:188] ^ 0);
  assign w706[31] = |(datain[187:184] ^ 0);
  assign w706[32] = |(datain[183:180] ^ 4);
  assign w706[33] = |(datain[179:176] ^ 2);
  assign w706[34] = |(datain[175:172] ^ 12);
  assign w706[35] = |(datain[171:168] ^ 13);
  assign w706[36] = |(datain[167:164] ^ 2);
  assign w706[37] = |(datain[163:160] ^ 1);
  assign w706[38] = |(datain[159:156] ^ 11);
  assign w706[39] = |(datain[155:152] ^ 4);
  assign w706[40] = |(datain[151:148] ^ 4);
  assign w706[41] = |(datain[147:144] ^ 0);
  assign w706[42] = |(datain[143:140] ^ 11);
  assign w706[43] = |(datain[139:136] ^ 10);
  assign w706[44] = |(datain[135:132] ^ 12);
  assign w706[45] = |(datain[131:128] ^ 2);
  assign comp[706] = ~(|w706);
  wire [46-1:0] w707;
  assign w707[0] = |(datain[311:308] ^ 13);
  assign w707[1] = |(datain[307:304] ^ 8);
  assign w707[2] = |(datain[303:300] ^ 11);
  assign w707[3] = |(datain[299:296] ^ 4);
  assign w707[4] = |(datain[295:292] ^ 4);
  assign w707[5] = |(datain[291:288] ^ 0);
  assign w707[6] = |(datain[287:284] ^ 3);
  assign w707[7] = |(datain[283:280] ^ 3);
  assign w707[8] = |(datain[279:276] ^ 13);
  assign w707[9] = |(datain[275:272] ^ 2);
  assign w707[10] = |(datain[271:268] ^ 11);
  assign w707[11] = |(datain[267:264] ^ 9);
  assign w707[12] = |(datain[263:260] ^ 11);
  assign w707[13] = |(datain[259:256] ^ 12);
  assign w707[14] = |(datain[255:252] ^ 0);
  assign w707[15] = |(datain[251:248] ^ 2);
  assign w707[16] = |(datain[247:244] ^ 12);
  assign w707[17] = |(datain[243:240] ^ 13);
  assign w707[18] = |(datain[239:236] ^ 2);
  assign w707[19] = |(datain[235:232] ^ 1);
  assign w707[20] = |(datain[231:228] ^ 3);
  assign w707[21] = |(datain[227:224] ^ 3);
  assign w707[22] = |(datain[223:220] ^ 12);
  assign w707[23] = |(datain[219:216] ^ 9);
  assign w707[24] = |(datain[215:212] ^ 3);
  assign w707[25] = |(datain[211:208] ^ 3);
  assign w707[26] = |(datain[207:204] ^ 13);
  assign w707[27] = |(datain[203:200] ^ 2);
  assign w707[28] = |(datain[199:196] ^ 11);
  assign w707[29] = |(datain[195:192] ^ 8);
  assign w707[30] = |(datain[191:188] ^ 0);
  assign w707[31] = |(datain[187:184] ^ 0);
  assign w707[32] = |(datain[183:180] ^ 4);
  assign w707[33] = |(datain[179:176] ^ 2);
  assign w707[34] = |(datain[175:172] ^ 12);
  assign w707[35] = |(datain[171:168] ^ 13);
  assign w707[36] = |(datain[167:164] ^ 2);
  assign w707[37] = |(datain[163:160] ^ 1);
  assign w707[38] = |(datain[159:156] ^ 11);
  assign w707[39] = |(datain[155:152] ^ 4);
  assign w707[40] = |(datain[151:148] ^ 4);
  assign w707[41] = |(datain[147:144] ^ 0);
  assign w707[42] = |(datain[143:140] ^ 11);
  assign w707[43] = |(datain[139:136] ^ 10);
  assign w707[44] = |(datain[135:132] ^ 10);
  assign w707[45] = |(datain[131:128] ^ 7);
  assign comp[707] = ~(|w707);
  wire [46-1:0] w708;
  assign w708[0] = |(datain[311:308] ^ 2);
  assign w708[1] = |(datain[307:304] ^ 12);
  assign w708[2] = |(datain[303:300] ^ 11);
  assign w708[3] = |(datain[299:296] ^ 11);
  assign w708[4] = |(datain[295:292] ^ 11);
  assign w708[5] = |(datain[291:288] ^ 0);
  assign w708[6] = |(datain[287:284] ^ 11);
  assign w708[7] = |(datain[283:280] ^ 0);
  assign w708[8] = |(datain[279:276] ^ 11);
  assign w708[9] = |(datain[275:272] ^ 9);
  assign w708[10] = |(datain[271:268] ^ 11);
  assign w708[11] = |(datain[267:264] ^ 14);
  assign w708[12] = |(datain[263:260] ^ 11);
  assign w708[13] = |(datain[259:256] ^ 10);
  assign w708[14] = |(datain[255:252] ^ 12);
  assign w708[15] = |(datain[251:248] ^ 13);
  assign w708[16] = |(datain[247:244] ^ 2);
  assign w708[17] = |(datain[243:240] ^ 1);
  assign w708[18] = |(datain[239:236] ^ 8);
  assign w708[19] = |(datain[235:232] ^ 1);
  assign w708[20] = |(datain[231:228] ^ 15);
  assign w708[21] = |(datain[227:224] ^ 11);
  assign w708[22] = |(datain[223:220] ^ 11);
  assign w708[23] = |(datain[219:216] ^ 14);
  assign w708[24] = |(datain[215:212] ^ 11);
  assign w708[25] = |(datain[211:208] ^ 10);
  assign w708[26] = |(datain[207:204] ^ 7);
  assign w708[27] = |(datain[203:200] ^ 5);
  assign w708[28] = |(datain[199:196] ^ 4);
  assign w708[29] = |(datain[195:192] ^ 11);
  assign w708[30] = |(datain[191:188] ^ 8);
  assign w708[31] = |(datain[187:184] ^ 1);
  assign w708[32] = |(datain[183:180] ^ 15);
  assign w708[33] = |(datain[179:176] ^ 9);
  assign w708[34] = |(datain[175:172] ^ 11);
  assign w708[35] = |(datain[171:168] ^ 0);
  assign w708[36] = |(datain[167:164] ^ 11);
  assign w708[37] = |(datain[163:160] ^ 0);
  assign w708[38] = |(datain[159:156] ^ 7);
  assign w708[39] = |(datain[155:152] ^ 5);
  assign w708[40] = |(datain[151:148] ^ 4);
  assign w708[41] = |(datain[147:144] ^ 5);
  assign w708[42] = |(datain[143:140] ^ 2);
  assign w708[43] = |(datain[139:136] ^ 14);
  assign w708[44] = |(datain[135:132] ^ 8);
  assign w708[45] = |(datain[131:128] ^ 3);
  assign comp[708] = ~(|w708);
  wire [42-1:0] w709;
  assign w709[0] = |(datain[311:308] ^ 0);
  assign w709[1] = |(datain[307:304] ^ 1);
  assign w709[2] = |(datain[303:300] ^ 8);
  assign w709[3] = |(datain[299:296] ^ 11);
  assign w709[4] = |(datain[295:292] ^ 1);
  assign w709[5] = |(datain[291:288] ^ 6);
  assign w709[6] = |(datain[287:284] ^ 8);
  assign w709[7] = |(datain[283:280] ^ 10);
  assign w709[8] = |(datain[279:276] ^ 0);
  assign w709[9] = |(datain[275:272] ^ 1);
  assign w709[10] = |(datain[271:268] ^ 14);
  assign w709[11] = |(datain[267:264] ^ 8);
  assign w709[12] = |(datain[263:260] ^ 6);
  assign w709[13] = |(datain[259:256] ^ 2);
  assign w709[14] = |(datain[255:252] ^ 0);
  assign w709[15] = |(datain[251:248] ^ 0);
  assign w709[16] = |(datain[247:244] ^ 8);
  assign w709[17] = |(datain[243:240] ^ 8);
  assign w709[18] = |(datain[239:236] ^ 13);
  assign w709[19] = |(datain[235:232] ^ 15);
  assign w709[20] = |(datain[231:228] ^ 11);
  assign w709[21] = |(datain[227:224] ^ 4);
  assign w709[22] = |(datain[223:220] ^ 0);
  assign w709[23] = |(datain[219:216] ^ 3);
  assign w709[24] = |(datain[215:212] ^ 11);
  assign w709[25] = |(datain[211:208] ^ 0);
  assign w709[26] = |(datain[207:204] ^ 0);
  assign w709[27] = |(datain[203:200] ^ 9);
  assign w709[28] = |(datain[199:196] ^ 14);
  assign w709[29] = |(datain[195:192] ^ 8);
  assign w709[30] = |(datain[191:188] ^ 5);
  assign w709[31] = |(datain[187:184] ^ 9);
  assign w709[32] = |(datain[183:180] ^ 0);
  assign w709[33] = |(datain[179:176] ^ 0);
  assign w709[34] = |(datain[175:172] ^ 11);
  assign w709[35] = |(datain[171:168] ^ 4);
  assign w709[36] = |(datain[167:164] ^ 0);
  assign w709[37] = |(datain[163:160] ^ 3);
  assign w709[38] = |(datain[159:156] ^ 11);
  assign w709[39] = |(datain[155:152] ^ 0);
  assign w709[40] = |(datain[151:148] ^ 0);
  assign w709[41] = |(datain[147:144] ^ 1);
  assign comp[709] = ~(|w709);
  wire [44-1:0] w710;
  assign w710[0] = |(datain[311:308] ^ 2);
  assign w710[1] = |(datain[307:304] ^ 6);
  assign w710[2] = |(datain[303:300] ^ 8);
  assign w710[3] = |(datain[299:296] ^ 8);
  assign w710[4] = |(datain[295:292] ^ 6);
  assign w710[5] = |(datain[291:288] ^ 5);
  assign w710[6] = |(datain[287:284] ^ 15);
  assign w710[7] = |(datain[283:280] ^ 14);
  assign w710[8] = |(datain[279:276] ^ 5);
  assign w710[9] = |(datain[275:272] ^ 15);
  assign w710[10] = |(datain[271:268] ^ 12);
  assign w710[11] = |(datain[267:264] ^ 13);
  assign w710[12] = |(datain[263:260] ^ 2);
  assign w710[13] = |(datain[259:256] ^ 1);
  assign w710[14] = |(datain[255:252] ^ 11);
  assign w710[15] = |(datain[251:248] ^ 4);
  assign w710[16] = |(datain[247:244] ^ 3);
  assign w710[17] = |(datain[243:240] ^ 12);
  assign w710[18] = |(datain[239:236] ^ 11);
  assign w710[19] = |(datain[235:232] ^ 1);
  assign w710[20] = |(datain[231:228] ^ 0);
  assign w710[21] = |(datain[227:224] ^ 2);
  assign w710[22] = |(datain[223:220] ^ 12);
  assign w710[23] = |(datain[219:216] ^ 13);
  assign w710[24] = |(datain[215:212] ^ 2);
  assign w710[25] = |(datain[211:208] ^ 1);
  assign w710[26] = |(datain[207:204] ^ 0);
  assign w710[27] = |(datain[203:200] ^ 14);
  assign w710[28] = |(datain[199:196] ^ 1);
  assign w710[29] = |(datain[195:192] ^ 15);
  assign w710[30] = |(datain[191:188] ^ 9);
  assign w710[31] = |(datain[187:184] ^ 3);
  assign w710[32] = |(datain[183:180] ^ 11);
  assign w710[33] = |(datain[179:176] ^ 4);
  assign w710[34] = |(datain[175:172] ^ 4);
  assign w710[35] = |(datain[171:168] ^ 0);
  assign w710[36] = |(datain[167:164] ^ 11);
  assign w710[37] = |(datain[163:160] ^ 10);
  assign w710[38] = |(datain[159:156] ^ 0);
  assign w710[39] = |(datain[155:152] ^ 0);
  assign w710[40] = |(datain[151:148] ^ 0);
  assign w710[41] = |(datain[147:144] ^ 1);
  assign w710[42] = |(datain[143:140] ^ 12);
  assign w710[43] = |(datain[139:136] ^ 13);
  assign comp[710] = ~(|w710);
  wire [74-1:0] w711;
  assign w711[0] = |(datain[311:308] ^ 12);
  assign w711[1] = |(datain[307:304] ^ 13);
  assign w711[2] = |(datain[303:300] ^ 2);
  assign w711[3] = |(datain[299:296] ^ 1);
  assign w711[4] = |(datain[295:292] ^ 0);
  assign w711[5] = |(datain[291:288] ^ 6);
  assign w711[6] = |(datain[287:284] ^ 11);
  assign w711[7] = |(datain[283:280] ^ 4);
  assign w711[8] = |(datain[279:276] ^ 4);
  assign w711[9] = |(datain[275:272] ^ 10);
  assign w711[10] = |(datain[271:268] ^ 11);
  assign w711[11] = |(datain[267:264] ^ 11);
  assign w711[12] = |(datain[263:260] ^ 15);
  assign w711[13] = |(datain[259:256] ^ 15);
  assign w711[14] = |(datain[255:252] ^ 15);
  assign w711[15] = |(datain[251:248] ^ 15);
  assign w711[16] = |(datain[247:244] ^ 12);
  assign w711[17] = |(datain[243:240] ^ 13);
  assign w711[18] = |(datain[239:236] ^ 2);
  assign w711[19] = |(datain[235:232] ^ 1);
  assign w711[20] = |(datain[231:228] ^ 11);
  assign w711[21] = |(datain[227:224] ^ 4);
  assign w711[22] = |(datain[223:220] ^ 4);
  assign w711[23] = |(datain[219:216] ^ 10);
  assign w711[24] = |(datain[215:212] ^ 11);
  assign w711[25] = |(datain[211:208] ^ 10);
  assign w711[26] = |(datain[207:204] ^ 1);
  assign w711[27] = |(datain[203:200] ^ 8);
  assign w711[28] = |(datain[199:196] ^ 0);
  assign w711[29] = |(datain[195:192] ^ 0);
  assign w711[30] = |(datain[191:188] ^ 2);
  assign w711[31] = |(datain[187:184] ^ 6);
  assign w711[32] = |(datain[183:180] ^ 2);
  assign w711[33] = |(datain[179:176] ^ 9);
  assign w711[34] = |(datain[175:172] ^ 1);
  assign w711[35] = |(datain[171:168] ^ 6);
  assign w711[36] = |(datain[167:164] ^ 0);
  assign w711[37] = |(datain[163:160] ^ 2);
  assign w711[38] = |(datain[159:156] ^ 0);
  assign w711[39] = |(datain[155:152] ^ 0);
  assign w711[40] = |(datain[151:148] ^ 2);
  assign w711[41] = |(datain[147:144] ^ 11);
  assign w711[42] = |(datain[143:140] ^ 13);
  assign w711[43] = |(datain[139:136] ^ 10);
  assign w711[44] = |(datain[135:132] ^ 12);
  assign w711[45] = |(datain[131:128] ^ 13);
  assign w711[46] = |(datain[127:124] ^ 2);
  assign w711[47] = |(datain[123:120] ^ 1);
  assign w711[48] = |(datain[119:116] ^ 11);
  assign w711[49] = |(datain[115:112] ^ 4);
  assign w711[50] = |(datain[111:108] ^ 4);
  assign w711[51] = |(datain[107:104] ^ 8);
  assign w711[52] = |(datain[103:100] ^ 8);
  assign w711[53] = |(datain[99:96] ^ 11);
  assign w711[54] = |(datain[95:92] ^ 13);
  assign w711[55] = |(datain[91:88] ^ 10);
  assign w711[56] = |(datain[87:84] ^ 4);
  assign w711[57] = |(datain[83:80] ^ 11);
  assign w711[58] = |(datain[79:76] ^ 12);
  assign w711[59] = |(datain[75:72] ^ 13);
  assign w711[60] = |(datain[71:68] ^ 2);
  assign w711[61] = |(datain[67:64] ^ 1);
  assign w711[62] = |(datain[63:60] ^ 4);
  assign w711[63] = |(datain[59:56] ^ 8);
  assign w711[64] = |(datain[55:52] ^ 8);
  assign w711[65] = |(datain[51:48] ^ 14);
  assign w711[66] = |(datain[47:44] ^ 12);
  assign w711[67] = |(datain[43:40] ^ 0);
  assign w711[68] = |(datain[39:36] ^ 4);
  assign w711[69] = |(datain[35:32] ^ 0);
  assign w711[70] = |(datain[31:28] ^ 2);
  assign w711[71] = |(datain[27:24] ^ 6);
  assign w711[72] = |(datain[23:20] ^ 12);
  assign w711[73] = |(datain[19:16] ^ 7);
  assign comp[711] = ~(|w711);
  wire [44-1:0] w712;
  assign w712[0] = |(datain[311:308] ^ 0);
  assign w712[1] = |(datain[307:304] ^ 3);
  assign w712[2] = |(datain[303:300] ^ 13);
  assign w712[3] = |(datain[299:296] ^ 1);
  assign w712[4] = |(datain[295:292] ^ 14);
  assign w712[5] = |(datain[291:288] ^ 9);
  assign w712[6] = |(datain[287:284] ^ 8);
  assign w712[7] = |(datain[283:280] ^ 3);
  assign w712[8] = |(datain[279:276] ^ 14);
  assign w712[9] = |(datain[275:272] ^ 9);
  assign w712[10] = |(datain[271:268] ^ 1);
  assign w712[11] = |(datain[267:264] ^ 0);
  assign w712[12] = |(datain[263:260] ^ 2);
  assign w712[13] = |(datain[259:256] ^ 14);
  assign w712[14] = |(datain[255:252] ^ 3);
  assign w712[15] = |(datain[251:248] ^ 1);
  assign w712[16] = |(datain[247:244] ^ 0);
  assign w712[17] = |(datain[243:240] ^ 7);
  assign w712[18] = |(datain[239:236] ^ 8);
  assign w712[19] = |(datain[235:232] ^ 3);
  assign w712[20] = |(datain[231:228] ^ 12);
  assign w712[21] = |(datain[227:224] ^ 3);
  assign w712[22] = |(datain[223:220] ^ 0);
  assign w712[23] = |(datain[219:216] ^ 2);
  assign w712[24] = |(datain[215:212] ^ 14);
  assign w712[25] = |(datain[211:208] ^ 2);
  assign w712[26] = |(datain[207:204] ^ 15);
  assign w712[27] = |(datain[203:200] ^ 8);
  assign w712[28] = |(datain[199:196] ^ 12);
  assign w712[29] = |(datain[195:192] ^ 3);
  assign w712[30] = |(datain[191:188] ^ 2);
  assign w712[31] = |(datain[187:184] ^ 14);
  assign w712[32] = |(datain[183:180] ^ 10);
  assign w712[33] = |(datain[179:176] ^ 3);
  assign w712[34] = |(datain[175:172] ^ 13);
  assign w712[35] = |(datain[171:168] ^ 8);
  assign w712[36] = |(datain[167:164] ^ 0);
  assign w712[37] = |(datain[163:160] ^ 14);
  assign w712[38] = |(datain[159:156] ^ 2);
  assign w712[39] = |(datain[155:152] ^ 14);
  assign w712[40] = |(datain[151:148] ^ 8);
  assign w712[41] = |(datain[147:144] ^ 9);
  assign w712[42] = |(datain[143:140] ^ 1);
  assign w712[43] = |(datain[139:136] ^ 14);
  assign comp[712] = ~(|w712);
  wire [40-1:0] w713;
  assign w713[0] = |(datain[311:308] ^ 14);
  assign w713[1] = |(datain[307:304] ^ 9);
  assign w713[2] = |(datain[303:300] ^ 8);
  assign w713[3] = |(datain[299:296] ^ 3);
  assign w713[4] = |(datain[295:292] ^ 14);
  assign w713[5] = |(datain[291:288] ^ 9);
  assign w713[6] = |(datain[287:284] ^ 1);
  assign w713[7] = |(datain[283:280] ^ 0);
  assign w713[8] = |(datain[279:276] ^ 2);
  assign w713[9] = |(datain[275:272] ^ 14);
  assign w713[10] = |(datain[271:268] ^ 3);
  assign w713[11] = |(datain[267:264] ^ 1);
  assign w713[12] = |(datain[263:260] ^ 0);
  assign w713[13] = |(datain[259:256] ^ 7);
  assign w713[14] = |(datain[255:252] ^ 8);
  assign w713[15] = |(datain[251:248] ^ 3);
  assign w713[16] = |(datain[247:244] ^ 12);
  assign w713[17] = |(datain[243:240] ^ 3);
  assign w713[18] = |(datain[239:236] ^ 0);
  assign w713[19] = |(datain[235:232] ^ 2);
  assign w713[20] = |(datain[231:228] ^ 14);
  assign w713[21] = |(datain[227:224] ^ 2);
  assign w713[22] = |(datain[223:220] ^ 15);
  assign w713[23] = |(datain[219:216] ^ 8);
  assign w713[24] = |(datain[215:212] ^ 12);
  assign w713[25] = |(datain[211:208] ^ 3);
  assign w713[26] = |(datain[207:204] ^ 2);
  assign w713[27] = |(datain[203:200] ^ 14);
  assign w713[28] = |(datain[199:196] ^ 10);
  assign w713[29] = |(datain[195:192] ^ 3);
  assign w713[30] = |(datain[191:188] ^ 6);
  assign w713[31] = |(datain[187:184] ^ 8);
  assign w713[32] = |(datain[183:180] ^ 0);
  assign w713[33] = |(datain[179:176] ^ 15);
  assign w713[34] = |(datain[175:172] ^ 2);
  assign w713[35] = |(datain[171:168] ^ 14);
  assign w713[36] = |(datain[167:164] ^ 8);
  assign w713[37] = |(datain[163:160] ^ 9);
  assign w713[38] = |(datain[159:156] ^ 1);
  assign w713[39] = |(datain[155:152] ^ 14);
  assign comp[713] = ~(|w713);
  wire [46-1:0] w714;
  assign w714[0] = |(datain[311:308] ^ 9);
  assign w714[1] = |(datain[307:304] ^ 0);
  assign w714[2] = |(datain[303:300] ^ 3);
  assign w714[3] = |(datain[299:296] ^ 3);
  assign w714[4] = |(datain[295:292] ^ 13);
  assign w714[5] = |(datain[291:288] ^ 9);
  assign w714[6] = |(datain[287:284] ^ 5);
  assign w714[7] = |(datain[283:280] ^ 3);
  assign w714[8] = |(datain[279:276] ^ 8);
  assign w714[9] = |(datain[275:272] ^ 11);
  assign w714[10] = |(datain[271:268] ^ 13);
  assign w714[11] = |(datain[267:264] ^ 5);
  assign w714[12] = |(datain[263:260] ^ 8);
  assign w714[13] = |(datain[259:256] ^ 3);
  assign w714[14] = |(datain[255:252] ^ 12);
  assign w714[15] = |(datain[251:248] ^ 4);
  assign w714[16] = |(datain[247:244] ^ 0);
  assign w714[17] = |(datain[243:240] ^ 2);
  assign w714[18] = |(datain[239:236] ^ 8);
  assign w714[19] = |(datain[235:232] ^ 11);
  assign w714[20] = |(datain[231:228] ^ 14);
  assign w714[21] = |(datain[227:224] ^ 12);
  assign w714[22] = |(datain[223:220] ^ 8);
  assign w714[23] = |(datain[219:216] ^ 3);
  assign w714[24] = |(datain[215:212] ^ 14);
  assign w714[25] = |(datain[211:208] ^ 13);
  assign w714[26] = |(datain[207:204] ^ 0);
  assign w714[27] = |(datain[203:200] ^ 2);
  assign w714[28] = |(datain[199:196] ^ 3);
  assign w714[29] = |(datain[195:192] ^ 1);
  assign w714[30] = |(datain[191:188] ^ 4);
  assign w714[31] = |(datain[187:184] ^ 14);
  assign w714[32] = |(datain[183:180] ^ 0);
  assign w714[33] = |(datain[179:176] ^ 0);
  assign w714[34] = |(datain[175:172] ^ 8);
  assign w714[35] = |(datain[171:168] ^ 3);
  assign w714[36] = |(datain[167:164] ^ 14);
  assign w714[37] = |(datain[163:160] ^ 12);
  assign w714[38] = |(datain[159:156] ^ 0);
  assign w714[39] = |(datain[155:152] ^ 2);
  assign w714[40] = |(datain[151:148] ^ 8);
  assign w714[41] = |(datain[147:144] ^ 11);
  assign w714[42] = |(datain[143:140] ^ 14);
  assign w714[43] = |(datain[139:136] ^ 10);
  assign w714[44] = |(datain[135:132] ^ 12);
  assign w714[45] = |(datain[131:128] ^ 3);
  assign comp[714] = ~(|w714);
  wire [44-1:0] w715;
  assign w715[0] = |(datain[311:308] ^ 2);
  assign w715[1] = |(datain[307:304] ^ 6);
  assign w715[2] = |(datain[303:300] ^ 8);
  assign w715[3] = |(datain[299:296] ^ 0);
  assign w715[4] = |(datain[295:292] ^ 7);
  assign w715[5] = |(datain[291:288] ^ 12);
  assign w715[6] = |(datain[287:284] ^ 0);
  assign w715[7] = |(datain[283:280] ^ 1);
  assign w715[8] = |(datain[279:276] ^ 3);
  assign w715[9] = |(datain[275:272] ^ 10);
  assign w715[10] = |(datain[271:268] ^ 7);
  assign w715[11] = |(datain[267:264] ^ 5);
  assign w715[12] = |(datain[263:260] ^ 0);
  assign w715[13] = |(datain[259:256] ^ 6);
  assign w715[14] = |(datain[255:252] ^ 2);
  assign w715[15] = |(datain[251:248] ^ 6);
  assign w715[16] = |(datain[247:244] ^ 8);
  assign w715[17] = |(datain[243:240] ^ 10);
  assign w715[18] = |(datain[239:236] ^ 1);
  assign w715[19] = |(datain[235:232] ^ 4);
  assign w715[20] = |(datain[231:228] ^ 8);
  assign w715[21] = |(datain[227:224] ^ 0);
  assign w715[22] = |(datain[223:220] ^ 14);
  assign w715[23] = |(datain[219:216] ^ 10);
  assign w715[24] = |(datain[215:212] ^ 4);
  assign w715[25] = |(datain[211:208] ^ 0);
  assign w715[26] = |(datain[207:204] ^ 11);
  assign w715[27] = |(datain[203:200] ^ 4);
  assign w715[28] = |(datain[199:196] ^ 3);
  assign w715[29] = |(datain[195:192] ^ 6);
  assign w715[30] = |(datain[191:188] ^ 14);
  assign w715[31] = |(datain[187:184] ^ 8);
  assign w715[32] = |(datain[183:180] ^ 13);
  assign w715[33] = |(datain[179:176] ^ 14);
  assign w715[34] = |(datain[175:172] ^ 15);
  assign w715[35] = |(datain[171:168] ^ 15);
  assign w715[36] = |(datain[167:164] ^ 3);
  assign w715[37] = |(datain[163:160] ^ 13);
  assign w715[38] = |(datain[159:156] ^ 15);
  assign w715[39] = |(datain[155:152] ^ 15);
  assign w715[40] = |(datain[151:148] ^ 15);
  assign w715[41] = |(datain[147:144] ^ 15);
  assign w715[42] = |(datain[143:140] ^ 7);
  assign w715[43] = |(datain[139:136] ^ 4);
  assign comp[715] = ~(|w715);
  wire [42-1:0] w716;
  assign w716[0] = |(datain[311:308] ^ 2);
  assign w716[1] = |(datain[307:304] ^ 2);
  assign w716[2] = |(datain[303:300] ^ 12);
  assign w716[3] = |(datain[299:296] ^ 13);
  assign w716[4] = |(datain[295:292] ^ 1);
  assign w716[5] = |(datain[291:288] ^ 3);
  assign w716[6] = |(datain[287:284] ^ 7);
  assign w716[7] = |(datain[283:280] ^ 2);
  assign w716[8] = |(datain[279:276] ^ 0);
  assign w716[9] = |(datain[275:272] ^ 3);
  assign w716[10] = |(datain[271:268] ^ 14);
  assign w716[11] = |(datain[267:264] ^ 9);
  assign w716[12] = |(datain[263:260] ^ 7);
  assign w716[13] = |(datain[259:256] ^ 1);
  assign w716[14] = |(datain[255:252] ^ 0);
  assign w716[15] = |(datain[251:248] ^ 2);
  assign w716[16] = |(datain[247:244] ^ 12);
  assign w716[17] = |(datain[243:240] ^ 6);
  assign w716[18] = |(datain[239:236] ^ 0);
  assign w716[19] = |(datain[235:232] ^ 6);
  assign w716[20] = |(datain[231:228] ^ 1);
  assign w716[21] = |(datain[227:224] ^ 15);
  assign w716[22] = |(datain[223:220] ^ 0);
  assign w716[23] = |(datain[219:216] ^ 8);
  assign w716[24] = |(datain[215:212] ^ 0);
  assign w716[25] = |(datain[211:208] ^ 0);
  assign w716[26] = |(datain[207:204] ^ 0);
  assign w716[27] = |(datain[203:200] ^ 14);
  assign w716[28] = |(datain[199:196] ^ 1);
  assign w716[29] = |(datain[195:192] ^ 15);
  assign w716[30] = |(datain[191:188] ^ 11);
  assign w716[31] = |(datain[187:184] ^ 8);
  assign w716[32] = |(datain[183:180] ^ 0);
  assign w716[33] = |(datain[179:176] ^ 0);
  assign w716[34] = |(datain[175:172] ^ 3);
  assign w716[35] = |(datain[171:168] ^ 13);
  assign w716[36] = |(datain[167:164] ^ 11);
  assign w716[37] = |(datain[163:160] ^ 10);
  assign w716[38] = |(datain[159:156] ^ 2);
  assign w716[39] = |(datain[155:152] ^ 4);
  assign w716[40] = |(datain[151:148] ^ 0);
  assign w716[41] = |(datain[147:144] ^ 8);
  assign comp[716] = ~(|w716);
  wire [76-1:0] w717;
  assign w717[0] = |(datain[311:308] ^ 2);
  assign w717[1] = |(datain[307:304] ^ 8);
  assign w717[2] = |(datain[303:300] ^ 0);
  assign w717[3] = |(datain[299:296] ^ 8);
  assign w717[4] = |(datain[295:292] ^ 0);
  assign w717[5] = |(datain[291:288] ^ 0);
  assign w717[6] = |(datain[287:284] ^ 10);
  assign w717[7] = |(datain[283:280] ^ 1);
  assign w717[8] = |(datain[279:276] ^ 3);
  assign w717[9] = |(datain[275:272] ^ 10);
  assign w717[10] = |(datain[271:268] ^ 0);
  assign w717[11] = |(datain[267:264] ^ 4);
  assign w717[12] = |(datain[263:260] ^ 10);
  assign w717[13] = |(datain[259:256] ^ 3);
  assign w717[14] = |(datain[255:252] ^ 3);
  assign w717[15] = |(datain[251:248] ^ 4);
  assign w717[16] = |(datain[247:244] ^ 0);
  assign w717[17] = |(datain[243:240] ^ 4);
  assign w717[18] = |(datain[239:236] ^ 10);
  assign w717[19] = |(datain[235:232] ^ 1);
  assign w717[20] = |(datain[231:228] ^ 3);
  assign w717[21] = |(datain[227:224] ^ 12);
  assign w717[22] = |(datain[223:220] ^ 0);
  assign w717[23] = |(datain[219:216] ^ 4);
  assign w717[24] = |(datain[215:212] ^ 10);
  assign w717[25] = |(datain[211:208] ^ 3);
  assign w717[26] = |(datain[207:204] ^ 3);
  assign w717[27] = |(datain[203:200] ^ 6);
  assign w717[28] = |(datain[199:196] ^ 0);
  assign w717[29] = |(datain[195:192] ^ 4);
  assign w717[30] = |(datain[191:188] ^ 10);
  assign w717[31] = |(datain[187:184] ^ 1);
  assign w717[32] = |(datain[183:180] ^ 3);
  assign w717[33] = |(datain[179:176] ^ 14);
  assign w717[34] = |(datain[175:172] ^ 0);
  assign w717[35] = |(datain[171:168] ^ 4);
  assign w717[36] = |(datain[167:164] ^ 10);
  assign w717[37] = |(datain[163:160] ^ 3);
  assign w717[38] = |(datain[159:156] ^ 3);
  assign w717[39] = |(datain[155:152] ^ 8);
  assign w717[40] = |(datain[151:148] ^ 0);
  assign w717[41] = |(datain[147:144] ^ 4);
  assign w717[42] = |(datain[143:140] ^ 15);
  assign w717[43] = |(datain[139:136] ^ 8);
  assign w717[44] = |(datain[135:132] ^ 11);
  assign w717[45] = |(datain[131:128] ^ 8);
  assign w717[46] = |(datain[127:124] ^ 0);
  assign w717[47] = |(datain[123:120] ^ 0);
  assign w717[48] = |(datain[119:116] ^ 2);
  assign w717[49] = |(datain[115:112] ^ 2);
  assign w717[50] = |(datain[111:108] ^ 12);
  assign w717[51] = |(datain[107:104] ^ 13);
  assign w717[52] = |(datain[103:100] ^ 1);
  assign w717[53] = |(datain[99:96] ^ 3);
  assign w717[54] = |(datain[95:92] ^ 7);
  assign w717[55] = |(datain[91:88] ^ 2);
  assign w717[56] = |(datain[87:84] ^ 0);
  assign w717[57] = |(datain[83:80] ^ 3);
  assign w717[58] = |(datain[79:76] ^ 14);
  assign w717[59] = |(datain[75:72] ^ 9);
  assign w717[60] = |(datain[71:68] ^ 7);
  assign w717[61] = |(datain[67:64] ^ 1);
  assign w717[62] = |(datain[63:60] ^ 0);
  assign w717[63] = |(datain[59:56] ^ 2);
  assign w717[64] = |(datain[55:52] ^ 12);
  assign w717[65] = |(datain[51:48] ^ 6);
  assign w717[66] = |(datain[47:44] ^ 0);
  assign w717[67] = |(datain[43:40] ^ 6);
  assign w717[68] = |(datain[39:36] ^ 2);
  assign w717[69] = |(datain[35:32] ^ 4);
  assign w717[70] = |(datain[31:28] ^ 0);
  assign w717[71] = |(datain[27:24] ^ 8);
  assign w717[72] = |(datain[23:20] ^ 0);
  assign w717[73] = |(datain[19:16] ^ 0);
  assign w717[74] = |(datain[15:12] ^ 0);
  assign w717[75] = |(datain[11:8] ^ 14);
  assign comp[717] = ~(|w717);
  wire [32-1:0] w718;
  assign w718[0] = |(datain[311:308] ^ 2);
  assign w718[1] = |(datain[307:304] ^ 1);
  assign w718[2] = |(datain[303:300] ^ 2);
  assign w718[3] = |(datain[299:296] ^ 5);
  assign w718[4] = |(datain[295:292] ^ 12);
  assign w718[5] = |(datain[291:288] ^ 13);
  assign w718[6] = |(datain[287:284] ^ 2);
  assign w718[7] = |(datain[283:280] ^ 1);
  assign w718[8] = |(datain[279:276] ^ 8);
  assign w718[9] = |(datain[275:272] ^ 12);
  assign w718[10] = |(datain[271:268] ^ 12);
  assign w718[11] = |(datain[267:264] ^ 8);
  assign w718[12] = |(datain[263:260] ^ 8);
  assign w718[13] = |(datain[259:256] ^ 14);
  assign w718[14] = |(datain[255:252] ^ 13);
  assign w718[15] = |(datain[251:248] ^ 8);
  assign w718[16] = |(datain[247:244] ^ 8);
  assign w718[17] = |(datain[243:240] ^ 14);
  assign w718[18] = |(datain[239:236] ^ 12);
  assign w718[19] = |(datain[235:232] ^ 0);
  assign w718[20] = |(datain[231:228] ^ 5);
  assign w718[21] = |(datain[227:224] ^ 8);
  assign w718[22] = |(datain[223:220] ^ 11);
  assign w718[23] = |(datain[219:216] ^ 11);
  assign w718[24] = |(datain[215:212] ^ 0);
  assign w718[25] = |(datain[211:208] ^ 0);
  assign w718[26] = |(datain[207:204] ^ 0);
  assign w718[27] = |(datain[203:200] ^ 1);
  assign w718[28] = |(datain[199:196] ^ 5);
  assign w718[29] = |(datain[195:192] ^ 3);
  assign w718[30] = |(datain[191:188] ^ 12);
  assign w718[31] = |(datain[187:184] ^ 3);
  assign comp[718] = ~(|w718);
  wire [30-1:0] w719;
  assign w719[0] = |(datain[311:308] ^ 2);
  assign w719[1] = |(datain[307:304] ^ 5);
  assign w719[2] = |(datain[303:300] ^ 12);
  assign w719[3] = |(datain[299:296] ^ 13);
  assign w719[4] = |(datain[295:292] ^ 2);
  assign w719[5] = |(datain[291:288] ^ 1);
  assign w719[6] = |(datain[287:284] ^ 8);
  assign w719[7] = |(datain[283:280] ^ 12);
  assign w719[8] = |(datain[279:276] ^ 12);
  assign w719[9] = |(datain[275:272] ^ 8);
  assign w719[10] = |(datain[271:268] ^ 8);
  assign w719[11] = |(datain[267:264] ^ 14);
  assign w719[12] = |(datain[263:260] ^ 13);
  assign w719[13] = |(datain[259:256] ^ 8);
  assign w719[14] = |(datain[255:252] ^ 8);
  assign w719[15] = |(datain[251:248] ^ 14);
  assign w719[16] = |(datain[247:244] ^ 12);
  assign w719[17] = |(datain[243:240] ^ 0);
  assign w719[18] = |(datain[239:236] ^ 5);
  assign w719[19] = |(datain[235:232] ^ 8);
  assign w719[20] = |(datain[231:228] ^ 11);
  assign w719[21] = |(datain[227:224] ^ 11);
  assign w719[22] = |(datain[223:220] ^ 0);
  assign w719[23] = |(datain[219:216] ^ 0);
  assign w719[24] = |(datain[215:212] ^ 0);
  assign w719[25] = |(datain[211:208] ^ 1);
  assign w719[26] = |(datain[207:204] ^ 5);
  assign w719[27] = |(datain[203:200] ^ 3);
  assign w719[28] = |(datain[199:196] ^ 12);
  assign w719[29] = |(datain[195:192] ^ 3);
  assign comp[719] = ~(|w719);
  wire [38-1:0] w720;
  assign w720[0] = |(datain[311:308] ^ 2);
  assign w720[1] = |(datain[307:304] ^ 1);
  assign w720[2] = |(datain[303:300] ^ 7);
  assign w720[3] = |(datain[299:296] ^ 2);
  assign w720[4] = |(datain[295:292] ^ 1);
  assign w720[5] = |(datain[291:288] ^ 9);
  assign w720[6] = |(datain[287:284] ^ 3);
  assign w720[7] = |(datain[283:280] ^ 11);
  assign w720[8] = |(datain[279:276] ^ 12);
  assign w720[9] = |(datain[275:272] ^ 1);
  assign w720[10] = |(datain[271:268] ^ 7);
  assign w720[11] = |(datain[267:264] ^ 2);
  assign w720[12] = |(datain[263:260] ^ 1);
  assign w720[13] = |(datain[259:256] ^ 5);
  assign w720[14] = |(datain[255:252] ^ 3);
  assign w720[15] = |(datain[251:248] ^ 3);
  assign w720[16] = |(datain[247:244] ^ 12);
  assign w720[17] = |(datain[243:240] ^ 9);
  assign w720[18] = |(datain[239:236] ^ 3);
  assign w720[19] = |(datain[235:232] ^ 3);
  assign w720[20] = |(datain[231:228] ^ 13);
  assign w720[21] = |(datain[227:224] ^ 2);
  assign w720[22] = |(datain[223:220] ^ 11);
  assign w720[23] = |(datain[219:216] ^ 8);
  assign w720[24] = |(datain[215:212] ^ 0);
  assign w720[25] = |(datain[211:208] ^ 0);
  assign w720[26] = |(datain[207:204] ^ 4);
  assign w720[27] = |(datain[203:200] ^ 2);
  assign w720[28] = |(datain[199:196] ^ 12);
  assign w720[29] = |(datain[195:192] ^ 13);
  assign w720[30] = |(datain[191:188] ^ 2);
  assign w720[31] = |(datain[187:184] ^ 1);
  assign w720[32] = |(datain[183:180] ^ 7);
  assign w720[33] = |(datain[179:176] ^ 2);
  assign w720[34] = |(datain[175:172] ^ 0);
  assign w720[35] = |(datain[171:168] ^ 10);
  assign w720[36] = |(datain[167:164] ^ 11);
  assign w720[37] = |(datain[163:160] ^ 10);
  assign comp[720] = ~(|w720);
  wire [44-1:0] w721;
  assign w721[0] = |(datain[311:308] ^ 0);
  assign w721[1] = |(datain[307:304] ^ 1);
  assign w721[2] = |(datain[303:300] ^ 8);
  assign w721[3] = |(datain[299:296] ^ 11);
  assign w721[4] = |(datain[295:292] ^ 1);
  assign w721[5] = |(datain[291:288] ^ 15);
  assign w721[6] = |(datain[287:284] ^ 11);
  assign w721[7] = |(datain[283:280] ^ 14);
  assign w721[8] = |(datain[279:276] ^ 1);
  assign w721[9] = |(datain[275:272] ^ 15);
  assign w721[10] = |(datain[271:268] ^ 0);
  assign w721[11] = |(datain[267:264] ^ 1);
  assign w721[12] = |(datain[263:260] ^ 0);
  assign w721[13] = |(datain[259:256] ^ 3);
  assign w721[14] = |(datain[255:252] ^ 15);
  assign w721[15] = |(datain[251:248] ^ 3);
  assign w721[16] = |(datain[247:244] ^ 11);
  assign w721[17] = |(datain[243:240] ^ 15);
  assign w721[18] = |(datain[239:236] ^ 0);
  assign w721[19] = |(datain[235:232] ^ 0);
  assign w721[20] = |(datain[231:228] ^ 0);
  assign w721[21] = |(datain[227:224] ^ 1);
  assign w721[22] = |(datain[223:220] ^ 11);
  assign w721[23] = |(datain[219:216] ^ 9);
  assign w721[24] = |(datain[215:212] ^ 0);
  assign w721[25] = |(datain[211:208] ^ 7);
  assign w721[26] = |(datain[207:204] ^ 0);
  assign w721[27] = |(datain[203:200] ^ 0);
  assign w721[28] = |(datain[199:196] ^ 15);
  assign w721[29] = |(datain[195:192] ^ 2);
  assign w721[30] = |(datain[191:188] ^ 10);
  assign w721[31] = |(datain[187:184] ^ 4);
  assign w721[32] = |(datain[183:180] ^ 14);
  assign w721[33] = |(datain[179:176] ^ 8);
  assign w721[34] = |(datain[175:172] ^ 0);
  assign w721[35] = |(datain[171:168] ^ 3);
  assign w721[36] = |(datain[167:164] ^ 0);
  assign w721[37] = |(datain[163:160] ^ 0);
  assign w721[38] = |(datain[159:156] ^ 0);
  assign w721[39] = |(datain[155:152] ^ 7);
  assign w721[40] = |(datain[151:148] ^ 1);
  assign w721[41] = |(datain[147:144] ^ 15);
  assign w721[42] = |(datain[143:140] ^ 12);
  assign w721[43] = |(datain[139:136] ^ 3);
  assign comp[721] = ~(|w721);
  wire [32-1:0] w722;
  assign w722[0] = |(datain[311:308] ^ 12);
  assign w722[1] = |(datain[307:304] ^ 3);
  assign w722[2] = |(datain[303:300] ^ 0);
  assign w722[3] = |(datain[299:296] ^ 2);
  assign w722[4] = |(datain[295:292] ^ 5);
  assign w722[5] = |(datain[291:288] ^ 3);
  assign w722[6] = |(datain[287:284] ^ 5);
  assign w722[7] = |(datain[283:280] ^ 1);
  assign w722[8] = |(datain[279:276] ^ 8);
  assign w722[9] = |(datain[275:272] ^ 11);
  assign w722[10] = |(datain[271:268] ^ 0);
  assign w722[11] = |(datain[267:264] ^ 7);
  assign w722[12] = |(datain[263:260] ^ 8);
  assign w722[13] = |(datain[259:256] ^ 11);
  assign w722[14] = |(datain[255:252] ^ 4);
  assign w722[15] = |(datain[251:248] ^ 15);
  assign w722[16] = |(datain[247:244] ^ 1);
  assign w722[17] = |(datain[243:240] ^ 0);
  assign w722[18] = |(datain[239:236] ^ 8);
  assign w722[19] = |(datain[235:232] ^ 11);
  assign w722[20] = |(datain[231:228] ^ 13);
  assign w722[21] = |(datain[227:224] ^ 8);
  assign w722[22] = |(datain[223:220] ^ 3);
  assign w722[23] = |(datain[219:216] ^ 0);
  assign w722[24] = |(datain[215:212] ^ 1);
  assign w722[25] = |(datain[211:208] ^ 15);
  assign w722[26] = |(datain[207:204] ^ 4);
  assign w722[27] = |(datain[203:200] ^ 3);
  assign w722[28] = |(datain[199:196] ^ 14);
  assign w722[29] = |(datain[195:192] ^ 2);
  assign w722[30] = |(datain[191:188] ^ 15);
  assign w722[31] = |(datain[187:184] ^ 11);
  assign comp[722] = ~(|w722);
  wire [76-1:0] w723;
  assign w723[0] = |(datain[311:308] ^ 12);
  assign w723[1] = |(datain[307:304] ^ 13);
  assign w723[2] = |(datain[303:300] ^ 2);
  assign w723[3] = |(datain[299:296] ^ 1);
  assign w723[4] = |(datain[295:292] ^ 11);
  assign w723[5] = |(datain[291:288] ^ 4);
  assign w723[6] = |(datain[287:284] ^ 1);
  assign w723[7] = |(datain[283:280] ^ 9);
  assign w723[8] = |(datain[279:276] ^ 12);
  assign w723[9] = |(datain[275:272] ^ 13);
  assign w723[10] = |(datain[271:268] ^ 2);
  assign w723[11] = |(datain[267:264] ^ 1);
  assign w723[12] = |(datain[263:260] ^ 8);
  assign w723[13] = |(datain[259:256] ^ 10);
  assign w723[14] = |(datain[255:252] ^ 13);
  assign w723[15] = |(datain[251:248] ^ 0);
  assign w723[16] = |(datain[247:244] ^ 15);
  assign w723[17] = |(datain[243:240] ^ 14);
  assign w723[18] = |(datain[239:236] ^ 12);
  assign w723[19] = |(datain[235:232] ^ 2);
  assign w723[20] = |(datain[231:228] ^ 11);
  assign w723[21] = |(datain[227:224] ^ 4);
  assign w723[22] = |(datain[223:220] ^ 4);
  assign w723[23] = |(datain[219:216] ^ 7);
  assign w723[24] = |(datain[215:212] ^ 11);
  assign w723[25] = |(datain[211:208] ^ 14);
  assign w723[26] = |(datain[207:204] ^ 4);
  assign w723[27] = |(datain[203:200] ^ 12);
  assign w723[28] = |(datain[199:196] ^ 0);
  assign w723[29] = |(datain[195:192] ^ 2);
  assign w723[30] = |(datain[191:188] ^ 12);
  assign w723[31] = |(datain[187:184] ^ 13);
  assign w723[32] = |(datain[183:180] ^ 2);
  assign w723[33] = |(datain[179:176] ^ 1);
  assign w723[34] = |(datain[175:172] ^ 11);
  assign w723[35] = |(datain[171:168] ^ 10);
  assign w723[36] = |(datain[167:164] ^ 14);
  assign w723[37] = |(datain[163:160] ^ 11);
  assign w723[38] = |(datain[159:156] ^ 0);
  assign w723[39] = |(datain[155:152] ^ 1);
  assign w723[40] = |(datain[151:148] ^ 11);
  assign w723[41] = |(datain[147:144] ^ 4);
  assign w723[42] = |(datain[143:140] ^ 3);
  assign w723[43] = |(datain[139:136] ^ 11);
  assign w723[44] = |(datain[135:132] ^ 12);
  assign w723[45] = |(datain[131:128] ^ 13);
  assign w723[46] = |(datain[127:124] ^ 2);
  assign w723[47] = |(datain[123:120] ^ 1);
  assign w723[48] = |(datain[119:116] ^ 11);
  assign w723[49] = |(datain[115:112] ^ 9);
  assign w723[50] = |(datain[111:108] ^ 1);
  assign w723[51] = |(datain[107:104] ^ 3);
  assign w723[52] = |(datain[103:100] ^ 0);
  assign w723[53] = |(datain[99:96] ^ 0);
  assign w723[54] = |(datain[95:92] ^ 11);
  assign w723[55] = |(datain[91:88] ^ 10);
  assign w723[56] = |(datain[87:84] ^ 14);
  assign w723[57] = |(datain[83:80] ^ 3);
  assign w723[58] = |(datain[79:76] ^ 0);
  assign w723[59] = |(datain[75:72] ^ 1);
  assign w723[60] = |(datain[71:68] ^ 11);
  assign w723[61] = |(datain[67:64] ^ 4);
  assign w723[62] = |(datain[63:60] ^ 4);
  assign w723[63] = |(datain[59:56] ^ 14);
  assign w723[64] = |(datain[55:52] ^ 12);
  assign w723[65] = |(datain[51:48] ^ 13);
  assign w723[66] = |(datain[47:44] ^ 2);
  assign w723[67] = |(datain[43:40] ^ 1);
  assign w723[68] = |(datain[39:36] ^ 3);
  assign w723[69] = |(datain[35:32] ^ 13);
  assign w723[70] = |(datain[31:28] ^ 1);
  assign w723[71] = |(datain[27:24] ^ 2);
  assign w723[72] = |(datain[23:20] ^ 0);
  assign w723[73] = |(datain[19:16] ^ 0);
  assign w723[74] = |(datain[15:12] ^ 7);
  assign w723[75] = |(datain[11:8] ^ 5);
  assign comp[723] = ~(|w723);
  wire [44-1:0] w724;
  assign w724[0] = |(datain[311:308] ^ 11);
  assign w724[1] = |(datain[307:304] ^ 10);
  assign w724[2] = |(datain[303:300] ^ 0);
  assign w724[3] = |(datain[299:296] ^ 0);
  assign w724[4] = |(datain[295:292] ^ 0);
  assign w724[5] = |(datain[291:288] ^ 1);
  assign w724[6] = |(datain[287:284] ^ 5);
  assign w724[7] = |(datain[283:280] ^ 9);
  assign w724[8] = |(datain[279:276] ^ 0);
  assign w724[9] = |(datain[275:272] ^ 3);
  assign w724[10] = |(datain[271:268] ^ 13);
  assign w724[11] = |(datain[267:264] ^ 1);
  assign w724[12] = |(datain[263:260] ^ 5);
  assign w724[13] = |(datain[259:256] ^ 1);
  assign w724[14] = |(datain[255:252] ^ 11);
  assign w724[15] = |(datain[251:248] ^ 9);
  assign w724[16] = |(datain[247:244] ^ 2);
  assign w724[17] = |(datain[243:240] ^ 13);
  assign w724[18] = |(datain[239:236] ^ 0);
  assign w724[19] = |(datain[235:232] ^ 2);
  assign w724[20] = |(datain[231:228] ^ 12);
  assign w724[21] = |(datain[227:224] ^ 13);
  assign w724[22] = |(datain[223:220] ^ 2);
  assign w724[23] = |(datain[219:216] ^ 1);
  assign w724[24] = |(datain[215:212] ^ 11);
  assign w724[25] = |(datain[211:208] ^ 15);
  assign w724[26] = |(datain[207:204] ^ 0);
  assign w724[27] = |(datain[203:200] ^ 1);
  assign w724[28] = |(datain[199:196] ^ 0);
  assign w724[29] = |(datain[195:192] ^ 3);
  assign w724[30] = |(datain[191:188] ^ 5);
  assign w724[31] = |(datain[187:184] ^ 9);
  assign w724[32] = |(datain[183:180] ^ 0);
  assign w724[33] = |(datain[179:176] ^ 3);
  assign w724[34] = |(datain[175:172] ^ 15);
  assign w724[35] = |(datain[171:168] ^ 9);
  assign w724[36] = |(datain[167:164] ^ 5);
  assign w724[37] = |(datain[163:160] ^ 1);
  assign w724[38] = |(datain[159:156] ^ 11);
  assign w724[39] = |(datain[155:152] ^ 9);
  assign w724[40] = |(datain[151:148] ^ 2);
  assign w724[41] = |(datain[147:144] ^ 6);
  assign w724[42] = |(datain[143:140] ^ 0);
  assign w724[43] = |(datain[139:136] ^ 0);
  assign comp[724] = ~(|w724);
  wire [42-1:0] w725;
  assign w725[0] = |(datain[311:308] ^ 0);
  assign w725[1] = |(datain[307:304] ^ 3);
  assign w725[2] = |(datain[303:300] ^ 15);
  assign w725[3] = |(datain[299:296] ^ 9);
  assign w725[4] = |(datain[295:292] ^ 11);
  assign w725[5] = |(datain[291:288] ^ 9);
  assign w725[6] = |(datain[287:284] ^ 2);
  assign w725[7] = |(datain[283:280] ^ 9);
  assign w725[8] = |(datain[279:276] ^ 0);
  assign w725[9] = |(datain[275:272] ^ 0);
  assign w725[10] = |(datain[271:268] ^ 3);
  assign w725[11] = |(datain[267:264] ^ 0);
  assign w725[12] = |(datain[263:260] ^ 3);
  assign w725[13] = |(datain[259:256] ^ 13);
  assign w725[14] = |(datain[255:252] ^ 4);
  assign w725[15] = |(datain[251:248] ^ 7);
  assign w725[16] = |(datain[247:244] ^ 14);
  assign w725[17] = |(datain[243:240] ^ 2);
  assign w725[18] = |(datain[239:236] ^ 15);
  assign w725[19] = |(datain[235:232] ^ 11);
  assign w725[20] = |(datain[231:228] ^ 15);
  assign w725[21] = |(datain[227:224] ^ 12);
  assign w725[22] = |(datain[223:220] ^ 11);
  assign w725[23] = |(datain[219:216] ^ 15);
  assign w725[24] = |(datain[215:212] ^ 0);
  assign w725[25] = |(datain[211:208] ^ 0);
  assign w725[26] = |(datain[207:204] ^ 0);
  assign w725[27] = |(datain[203:200] ^ 1);
  assign w725[28] = |(datain[199:196] ^ 11);
  assign w725[29] = |(datain[195:192] ^ 14);
  assign w725[30] = |(datain[191:188] ^ 3);
  assign w725[31] = |(datain[187:184] ^ 9);
  assign w725[32] = |(datain[183:180] ^ 0);
  assign w725[33] = |(datain[179:176] ^ 3);
  assign w725[34] = |(datain[175:172] ^ 5);
  assign w725[35] = |(datain[171:168] ^ 9);
  assign w725[36] = |(datain[167:164] ^ 0);
  assign w725[37] = |(datain[163:160] ^ 3);
  assign w725[38] = |(datain[159:156] ^ 15);
  assign w725[39] = |(datain[155:152] ^ 1);
  assign w725[40] = |(datain[151:148] ^ 5);
  assign w725[41] = |(datain[147:144] ^ 1);
  assign comp[725] = ~(|w725);
  wire [76-1:0] w726;
  assign w726[0] = |(datain[311:308] ^ 15);
  assign w726[1] = |(datain[307:304] ^ 7);
  assign w726[2] = |(datain[303:300] ^ 15);
  assign w726[3] = |(datain[299:296] ^ 1);
  assign w726[4] = |(datain[295:292] ^ 4);
  assign w726[5] = |(datain[291:288] ^ 0);
  assign w726[6] = |(datain[287:284] ^ 10);
  assign w726[7] = |(datain[283:280] ^ 3);
  assign w726[8] = |(datain[279:276] ^ 3);
  assign w726[9] = |(datain[275:272] ^ 8);
  assign w726[10] = |(datain[271:268] ^ 0);
  assign w726[11] = |(datain[267:264] ^ 1);
  assign w726[12] = |(datain[263:260] ^ 11);
  assign w726[13] = |(datain[259:256] ^ 4);
  assign w726[14] = |(datain[255:252] ^ 4);
  assign w726[15] = |(datain[251:248] ^ 0);
  assign w726[16] = |(datain[247:244] ^ 8);
  assign w726[17] = |(datain[243:240] ^ 11);
  assign w726[18] = |(datain[239:236] ^ 1);
  assign w726[19] = |(datain[235:232] ^ 14);
  assign w726[20] = |(datain[231:228] ^ 4);
  assign w726[21] = |(datain[227:224] ^ 0);
  assign w726[22] = |(datain[223:220] ^ 0);
  assign w726[23] = |(datain[219:216] ^ 1);
  assign w726[24] = |(datain[215:212] ^ 11);
  assign w726[25] = |(datain[211:208] ^ 9);
  assign w726[26] = |(datain[207:204] ^ 1);
  assign w726[27] = |(datain[203:200] ^ 0);
  assign w726[28] = |(datain[199:196] ^ 0);
  assign w726[29] = |(datain[195:192] ^ 0);
  assign w726[30] = |(datain[191:188] ^ 2);
  assign w726[31] = |(datain[187:184] ^ 9);
  assign w726[32] = |(datain[183:180] ^ 13);
  assign w726[33] = |(datain[179:176] ^ 1);
  assign w726[34] = |(datain[175:172] ^ 11);
  assign w726[35] = |(datain[171:168] ^ 10);
  assign w726[36] = |(datain[167:164] ^ 4);
  assign w726[37] = |(datain[163:160] ^ 4);
  assign w726[38] = |(datain[159:156] ^ 0);
  assign w726[39] = |(datain[155:152] ^ 1);
  assign w726[40] = |(datain[151:148] ^ 12);
  assign w726[41] = |(datain[147:144] ^ 13);
  assign w726[42] = |(datain[143:140] ^ 2);
  assign w726[43] = |(datain[139:136] ^ 1);
  assign w726[44] = |(datain[135:132] ^ 7);
  assign w726[45] = |(datain[131:128] ^ 2);
  assign w726[46] = |(datain[127:124] ^ 1);
  assign w726[47] = |(datain[123:120] ^ 15);
  assign w726[48] = |(datain[119:116] ^ 11);
  assign w726[49] = |(datain[115:112] ^ 8);
  assign w726[50] = |(datain[111:108] ^ 0);
  assign w726[51] = |(datain[107:104] ^ 0);
  assign w726[52] = |(datain[103:100] ^ 4);
  assign w726[53] = |(datain[99:96] ^ 2);
  assign w726[54] = |(datain[95:92] ^ 8);
  assign w726[55] = |(datain[91:88] ^ 11);
  assign w726[56] = |(datain[87:84] ^ 1);
  assign w726[57] = |(datain[83:80] ^ 14);
  assign w726[58] = |(datain[79:76] ^ 4);
  assign w726[59] = |(datain[75:72] ^ 0);
  assign w726[60] = |(datain[71:68] ^ 0);
  assign w726[61] = |(datain[67:64] ^ 1);
  assign w726[62] = |(datain[63:60] ^ 11);
  assign w726[63] = |(datain[59:56] ^ 9);
  assign w726[64] = |(datain[55:52] ^ 0);
  assign w726[65] = |(datain[51:48] ^ 0);
  assign w726[66] = |(datain[47:44] ^ 0);
  assign w726[67] = |(datain[43:40] ^ 0);
  assign w726[68] = |(datain[39:36] ^ 11);
  assign w726[69] = |(datain[35:32] ^ 10);
  assign w726[70] = |(datain[31:28] ^ 0);
  assign w726[71] = |(datain[27:24] ^ 0);
  assign w726[72] = |(datain[23:20] ^ 0);
  assign w726[73] = |(datain[19:16] ^ 0);
  assign w726[74] = |(datain[15:12] ^ 12);
  assign w726[75] = |(datain[11:8] ^ 13);
  assign comp[726] = ~(|w726);
  wire [68-1:0] w727;
  assign w727[0] = |(datain[311:308] ^ 5);
  assign w727[1] = |(datain[307:304] ^ 11);
  assign w727[2] = |(datain[303:300] ^ 8);
  assign w727[3] = |(datain[299:296] ^ 3);
  assign w727[4] = |(datain[295:292] ^ 14);
  assign w727[5] = |(datain[291:288] ^ 11);
  assign w727[6] = |(datain[287:284] ^ 0);
  assign w727[7] = |(datain[283:280] ^ 3);
  assign w727[8] = |(datain[279:276] ^ 15);
  assign w727[9] = |(datain[275:272] ^ 10);
  assign w727[10] = |(datain[271:268] ^ 8);
  assign w727[11] = |(datain[267:264] ^ 11);
  assign w727[12] = |(datain[263:260] ^ 12);
  assign w727[13] = |(datain[259:256] ^ 11);
  assign w727[14] = |(datain[255:252] ^ 8);
  assign w727[15] = |(datain[251:248] ^ 1);
  assign w727[16] = |(datain[247:244] ^ 14);
  assign w727[17] = |(datain[243:240] ^ 9);
  assign w727[18] = |(datain[239:236] ^ 0);
  assign w727[19] = |(datain[235:232] ^ 0);
  assign w727[20] = |(datain[231:228] ^ 0);
  assign w727[21] = |(datain[227:224] ^ 1);
  assign w727[22] = |(datain[223:220] ^ 8);
  assign w727[23] = |(datain[219:216] ^ 11);
  assign w727[24] = |(datain[215:212] ^ 14);
  assign w727[25] = |(datain[211:208] ^ 3);
  assign w727[26] = |(datain[207:204] ^ 8);
  assign w727[27] = |(datain[203:200] ^ 1);
  assign w727[28] = |(datain[199:196] ^ 12);
  assign w727[29] = |(datain[195:192] ^ 4);
  assign w727[30] = |(datain[191:188] ^ 2);
  assign w727[31] = |(datain[187:184] ^ 13);
  assign w727[32] = |(datain[183:180] ^ 0);
  assign w727[33] = |(datain[179:176] ^ 0);
  assign w727[34] = |(datain[175:172] ^ 5);
  assign w727[35] = |(datain[171:168] ^ 14);
  assign w727[36] = |(datain[167:164] ^ 8);
  assign w727[37] = |(datain[163:160] ^ 3);
  assign w727[38] = |(datain[159:156] ^ 14);
  assign w727[39] = |(datain[155:152] ^ 12);
  assign w727[40] = |(datain[151:148] ^ 0);
  assign w727[41] = |(datain[147:144] ^ 4);
  assign w727[42] = |(datain[143:140] ^ 5);
  assign w727[43] = |(datain[139:136] ^ 8);
  assign w727[44] = |(datain[135:132] ^ 8);
  assign w727[45] = |(datain[131:128] ^ 3);
  assign w727[46] = |(datain[127:124] ^ 14);
  assign w727[47] = |(datain[123:120] ^ 12);
  assign w727[48] = |(datain[119:116] ^ 0);
  assign w727[49] = |(datain[115:112] ^ 4);
  assign w727[50] = |(datain[111:108] ^ 15);
  assign w727[51] = |(datain[107:104] ^ 12);
  assign w727[52] = |(datain[103:100] ^ 3);
  assign w727[53] = |(datain[99:96] ^ 0);
  assign w727[54] = |(datain[95:92] ^ 0);
  assign w727[55] = |(datain[91:88] ^ 4);
  assign w727[56] = |(datain[87:84] ^ 4);
  assign w727[57] = |(datain[83:80] ^ 6);
  assign w727[58] = |(datain[79:76] ^ 14);
  assign w727[59] = |(datain[75:72] ^ 2);
  assign w727[60] = |(datain[71:68] ^ 15);
  assign w727[61] = |(datain[67:64] ^ 11);
  assign w727[62] = |(datain[63:60] ^ 14);
  assign w727[63] = |(datain[59:56] ^ 9);
  assign w727[64] = |(datain[55:52] ^ 7);
  assign w727[65] = |(datain[51:48] ^ 7);
  assign w727[66] = |(datain[47:44] ^ 15);
  assign w727[67] = |(datain[43:40] ^ 14);
  assign comp[727] = ~(|w727);
  wire [28-1:0] w728;
  assign w728[0] = |(datain[311:308] ^ 14);
  assign w728[1] = |(datain[307:304] ^ 11);
  assign w728[2] = |(datain[303:300] ^ 13);
  assign w728[3] = |(datain[299:296] ^ 9);
  assign w728[4] = |(datain[295:292] ^ 11);
  assign w728[5] = |(datain[291:288] ^ 4);
  assign w728[6] = |(datain[287:284] ^ 2);
  assign w728[7] = |(datain[283:280] ^ 10);
  assign w728[8] = |(datain[279:276] ^ 12);
  assign w728[9] = |(datain[275:272] ^ 13);
  assign w728[10] = |(datain[271:268] ^ 2);
  assign w728[11] = |(datain[267:264] ^ 1);
  assign w728[12] = |(datain[263:260] ^ 3);
  assign w728[13] = |(datain[259:256] ^ 12);
  assign w728[14] = |(datain[255:252] ^ 0);
  assign w728[15] = |(datain[251:248] ^ 1);
  assign w728[16] = |(datain[247:244] ^ 7);
  assign w728[17] = |(datain[243:240] ^ 4);
  assign w728[18] = |(datain[239:236] ^ 1);
  assign w728[19] = |(datain[235:232] ^ 1);
  assign w728[20] = |(datain[231:228] ^ 14);
  assign w728[21] = |(datain[227:224] ^ 11);
  assign w728[22] = |(datain[223:220] ^ 1);
  assign w728[23] = |(datain[219:216] ^ 13);
  assign w728[24] = |(datain[215:212] ^ 9);
  assign w728[25] = |(datain[211:208] ^ 0);
  assign w728[26] = |(datain[207:204] ^ 0);
  assign w728[27] = |(datain[203:200] ^ 7);
  assign comp[728] = ~(|w728);
  wire [30-1:0] w729;
  assign w729[0] = |(datain[311:308] ^ 14);
  assign w729[1] = |(datain[307:304] ^ 11);
  assign w729[2] = |(datain[303:300] ^ 13);
  assign w729[3] = |(datain[299:296] ^ 9);
  assign w729[4] = |(datain[295:292] ^ 11);
  assign w729[5] = |(datain[291:288] ^ 4);
  assign w729[6] = |(datain[287:284] ^ 2);
  assign w729[7] = |(datain[283:280] ^ 10);
  assign w729[8] = |(datain[279:276] ^ 12);
  assign w729[9] = |(datain[275:272] ^ 13);
  assign w729[10] = |(datain[271:268] ^ 2);
  assign w729[11] = |(datain[267:264] ^ 1);
  assign w729[12] = |(datain[263:260] ^ 3);
  assign w729[13] = |(datain[259:256] ^ 12);
  assign w729[14] = |(datain[255:252] ^ 0);
  assign w729[15] = |(datain[251:248] ^ 1);
  assign w729[16] = |(datain[247:244] ^ 7);
  assign w729[17] = |(datain[243:240] ^ 4);
  assign w729[18] = |(datain[239:236] ^ 1);
  assign w729[19] = |(datain[235:232] ^ 1);
  assign w729[20] = |(datain[231:228] ^ 14);
  assign w729[21] = |(datain[227:224] ^ 11);
  assign w729[22] = |(datain[223:220] ^ 1);
  assign w729[23] = |(datain[219:216] ^ 13);
  assign w729[24] = |(datain[215:212] ^ 9);
  assign w729[25] = |(datain[211:208] ^ 0);
  assign w729[26] = |(datain[207:204] ^ 0);
  assign w729[27] = |(datain[203:200] ^ 7);
  assign w729[28] = |(datain[199:196] ^ 1);
  assign w729[29] = |(datain[195:192] ^ 15);
  assign comp[729] = ~(|w729);
  wire [28-1:0] w730;
  assign w730[0] = |(datain[311:308] ^ 0);
  assign w730[1] = |(datain[307:304] ^ 1);
  assign w730[2] = |(datain[303:300] ^ 9);
  assign w730[3] = |(datain[299:296] ^ 0);
  assign w730[4] = |(datain[295:292] ^ 11);
  assign w730[5] = |(datain[291:288] ^ 9);
  assign w730[6] = |(datain[287:284] ^ 0);
  assign w730[7] = |(datain[283:280] ^ 11);
  assign w730[8] = |(datain[279:276] ^ 1);
  assign w730[9] = |(datain[275:272] ^ 1);
  assign w730[10] = |(datain[271:268] ^ 9);
  assign w730[11] = |(datain[267:264] ^ 0);
  assign w730[12] = |(datain[263:260] ^ 11);
  assign w730[13] = |(datain[259:256] ^ 4);
  assign w730[14] = |(datain[255:252] ^ 4);
  assign w730[15] = |(datain[251:248] ^ 14);
  assign w730[16] = |(datain[247:244] ^ 12);
  assign w730[17] = |(datain[243:240] ^ 13);
  assign w730[18] = |(datain[239:236] ^ 2);
  assign w730[19] = |(datain[235:232] ^ 1);
  assign w730[20] = |(datain[231:228] ^ 9);
  assign w730[21] = |(datain[227:224] ^ 0);
  assign w730[22] = |(datain[223:220] ^ 7);
  assign w730[23] = |(datain[219:216] ^ 3);
  assign w730[24] = |(datain[215:212] ^ 0);
  assign w730[25] = |(datain[211:208] ^ 3);
  assign w730[26] = |(datain[207:204] ^ 9);
  assign w730[27] = |(datain[203:200] ^ 0);
  assign comp[730] = ~(|w730);
  wire [28-1:0] w731;
  assign w731[0] = |(datain[311:308] ^ 0);
  assign w731[1] = |(datain[307:304] ^ 1);
  assign w731[2] = |(datain[303:300] ^ 11);
  assign w731[3] = |(datain[299:296] ^ 9);
  assign w731[4] = |(datain[295:292] ^ 0);
  assign w731[5] = |(datain[291:288] ^ 11);
  assign w731[6] = |(datain[287:284] ^ 1);
  assign w731[7] = |(datain[283:280] ^ 1);
  assign w731[8] = |(datain[279:276] ^ 9);
  assign w731[9] = |(datain[275:272] ^ 0);
  assign w731[10] = |(datain[271:268] ^ 11);
  assign w731[11] = |(datain[267:264] ^ 4);
  assign w731[12] = |(datain[263:260] ^ 4);
  assign w731[13] = |(datain[259:256] ^ 14);
  assign w731[14] = |(datain[255:252] ^ 12);
  assign w731[15] = |(datain[251:248] ^ 13);
  assign w731[16] = |(datain[247:244] ^ 2);
  assign w731[17] = |(datain[243:240] ^ 1);
  assign w731[18] = |(datain[239:236] ^ 9);
  assign w731[19] = |(datain[235:232] ^ 0);
  assign w731[20] = |(datain[231:228] ^ 7);
  assign w731[21] = |(datain[227:224] ^ 3);
  assign w731[22] = |(datain[223:220] ^ 0);
  assign w731[23] = |(datain[219:216] ^ 2);
  assign w731[24] = |(datain[215:212] ^ 14);
  assign w731[25] = |(datain[211:208] ^ 11);
  assign w731[26] = |(datain[207:204] ^ 2);
  assign w731[27] = |(datain[203:200] ^ 5);
  assign comp[731] = ~(|w731);
  wire [46-1:0] w732;
  assign w732[0] = |(datain[311:308] ^ 13);
  assign w732[1] = |(datain[307:304] ^ 8);
  assign w732[2] = |(datain[303:300] ^ 11);
  assign w732[3] = |(datain[299:296] ^ 14);
  assign w732[4] = |(datain[295:292] ^ 8);
  assign w732[5] = |(datain[291:288] ^ 4);
  assign w732[6] = |(datain[287:284] ^ 0);
  assign w732[7] = |(datain[283:280] ^ 0);
  assign w732[8] = |(datain[279:276] ^ 11);
  assign w732[9] = |(datain[275:272] ^ 15);
  assign w732[10] = |(datain[271:268] ^ 0);
  assign w732[11] = |(datain[267:264] ^ 14);
  assign w732[12] = |(datain[263:260] ^ 0);
  assign w732[13] = |(datain[259:256] ^ 0);
  assign w732[14] = |(datain[255:252] ^ 10);
  assign w732[15] = |(datain[251:248] ^ 5);
  assign w732[16] = |(datain[247:244] ^ 10);
  assign w732[17] = |(datain[243:240] ^ 5);
  assign w732[18] = |(datain[239:236] ^ 15);
  assign w732[19] = |(datain[235:232] ^ 10);
  assign w732[20] = |(datain[231:228] ^ 12);
  assign w732[21] = |(datain[227:224] ^ 7);
  assign w732[22] = |(datain[223:220] ^ 4);
  assign w732[23] = |(datain[219:216] ^ 4);
  assign w732[24] = |(datain[215:212] ^ 15);
  assign w732[25] = |(datain[211:208] ^ 12);
  assign w732[26] = |(datain[207:204] ^ 2);
  assign w732[27] = |(datain[203:200] ^ 10);
  assign w732[28] = |(datain[199:196] ^ 0);
  assign w732[29] = |(datain[195:192] ^ 0);
  assign w732[30] = |(datain[191:188] ^ 8);
  assign w732[31] = |(datain[187:184] ^ 12);
  assign w732[32] = |(datain[183:180] ^ 4);
  assign w732[33] = |(datain[179:176] ^ 4);
  assign w732[34] = |(datain[175:172] ^ 15);
  assign w732[35] = |(datain[171:168] ^ 14);
  assign w732[36] = |(datain[167:164] ^ 15);
  assign w732[37] = |(datain[163:160] ^ 11);
  assign w732[38] = |(datain[159:156] ^ 11);
  assign w732[39] = |(datain[155:152] ^ 14);
  assign w732[40] = |(datain[151:148] ^ 2);
  assign w732[41] = |(datain[147:144] ^ 0);
  assign w732[42] = |(datain[143:140] ^ 0);
  assign w732[43] = |(datain[139:136] ^ 0);
  assign w732[44] = |(datain[135:132] ^ 11);
  assign w732[45] = |(datain[131:128] ^ 15);
  assign comp[732] = ~(|w732);
  wire [76-1:0] w733;
  assign w733[0] = |(datain[311:308] ^ 0);
  assign w733[1] = |(datain[307:304] ^ 14);
  assign w733[2] = |(datain[303:300] ^ 4);
  assign w733[3] = |(datain[299:296] ^ 6);
  assign w733[4] = |(datain[295:292] ^ 0);
  assign w733[5] = |(datain[291:288] ^ 0);
  assign w733[6] = |(datain[287:284] ^ 14);
  assign w733[7] = |(datain[283:280] ^ 8);
  assign w733[8] = |(datain[279:276] ^ 1);
  assign w733[9] = |(datain[275:272] ^ 4);
  assign w733[10] = |(datain[271:268] ^ 0);
  assign w733[11] = |(datain[267:264] ^ 0);
  assign w733[12] = |(datain[263:260] ^ 5);
  assign w733[13] = |(datain[259:256] ^ 10);
  assign w733[14] = |(datain[255:252] ^ 5);
  assign w733[15] = |(datain[251:248] ^ 9);
  assign w733[16] = |(datain[247:244] ^ 7);
  assign w733[17] = |(datain[243:240] ^ 2);
  assign w733[18] = |(datain[239:236] ^ 0);
  assign w733[19] = |(datain[235:232] ^ 10);
  assign w733[20] = |(datain[231:228] ^ 14);
  assign w733[21] = |(datain[227:224] ^ 8);
  assign w733[22] = |(datain[223:220] ^ 3);
  assign w733[23] = |(datain[219:216] ^ 14);
  assign w733[24] = |(datain[215:212] ^ 15);
  assign w733[25] = |(datain[211:208] ^ 15);
  assign w733[26] = |(datain[207:204] ^ 3);
  assign w733[27] = |(datain[203:200] ^ 3);
  assign w733[28] = |(datain[199:196] ^ 13);
  assign w733[29] = |(datain[195:192] ^ 11);
  assign w733[30] = |(datain[191:188] ^ 14);
  assign w733[31] = |(datain[187:184] ^ 8);
  assign w733[32] = |(datain[183:180] ^ 0);
  assign w733[33] = |(datain[179:176] ^ 8);
  assign w733[34] = |(datain[175:172] ^ 0);
  assign w733[35] = |(datain[171:168] ^ 0);
  assign w733[36] = |(datain[167:164] ^ 3);
  assign w733[37] = |(datain[163:160] ^ 3);
  assign w733[38] = |(datain[159:156] ^ 15);
  assign w733[39] = |(datain[155:152] ^ 6);
  assign w733[40] = |(datain[151:148] ^ 5);
  assign w733[41] = |(datain[147:144] ^ 8);
  assign w733[42] = |(datain[143:140] ^ 5);
  assign w733[43] = |(datain[139:136] ^ 9);
  assign w733[44] = |(datain[135:132] ^ 5);
  assign w733[45] = |(datain[131:128] ^ 11);
  assign w733[46] = |(datain[127:124] ^ 1);
  assign w733[47] = |(datain[123:120] ^ 15);
  assign w733[48] = |(datain[119:116] ^ 0);
  assign w733[49] = |(datain[115:112] ^ 7);
  assign w733[50] = |(datain[111:108] ^ 12);
  assign w733[51] = |(datain[107:104] ^ 3);
  assign w733[52] = |(datain[103:100] ^ 11);
  assign w733[53] = |(datain[99:96] ^ 8);
  assign w733[54] = |(datain[95:92] ^ 0);
  assign w733[55] = |(datain[91:88] ^ 1);
  assign w733[56] = |(datain[87:84] ^ 0);
  assign w733[57] = |(datain[83:80] ^ 3);
  assign w733[58] = |(datain[79:76] ^ 14);
  assign w733[59] = |(datain[75:72] ^ 8);
  assign w733[60] = |(datain[71:68] ^ 1);
  assign w733[61] = |(datain[67:64] ^ 10);
  assign w733[62] = |(datain[63:60] ^ 15);
  assign w733[63] = |(datain[59:56] ^ 15);
  assign w733[64] = |(datain[55:52] ^ 12);
  assign w733[65] = |(datain[51:48] ^ 3);
  assign w733[66] = |(datain[47:44] ^ 8);
  assign w733[67] = |(datain[43:40] ^ 0);
  assign w733[68] = |(datain[39:36] ^ 15);
  assign w733[69] = |(datain[35:32] ^ 12);
  assign w733[70] = |(datain[31:28] ^ 0);
  assign w733[71] = |(datain[27:24] ^ 0);
  assign w733[72] = |(datain[23:20] ^ 7);
  assign w733[73] = |(datain[19:16] ^ 5);
  assign w733[74] = |(datain[15:12] ^ 0);
  assign w733[75] = |(datain[11:8] ^ 12);
  assign comp[733] = ~(|w733);
  wire [74-1:0] w734;
  assign w734[0] = |(datain[311:308] ^ 15);
  assign w734[1] = |(datain[307:304] ^ 2);
  assign w734[2] = |(datain[303:300] ^ 0);
  assign w734[3] = |(datain[299:296] ^ 2);
  assign w734[4] = |(datain[295:292] ^ 14);
  assign w734[5] = |(datain[291:288] ^ 8);
  assign w734[6] = |(datain[287:284] ^ 6);
  assign w734[7] = |(datain[283:280] ^ 9);
  assign w734[8] = |(datain[279:276] ^ 15);
  assign w734[9] = |(datain[275:272] ^ 15);
  assign w734[10] = |(datain[271:268] ^ 12);
  assign w734[11] = |(datain[267:264] ^ 3);
  assign w734[12] = |(datain[263:260] ^ 11);
  assign w734[13] = |(datain[259:256] ^ 4);
  assign w734[14] = |(datain[255:252] ^ 4);
  assign w734[15] = |(datain[251:248] ^ 3);
  assign w734[16] = |(datain[247:244] ^ 11);
  assign w734[17] = |(datain[243:240] ^ 0);
  assign w734[18] = |(datain[239:236] ^ 0);
  assign w734[19] = |(datain[235:232] ^ 1);
  assign w734[20] = |(datain[231:228] ^ 11);
  assign w734[21] = |(datain[227:224] ^ 10);
  assign w734[22] = |(datain[223:220] ^ 0);
  assign w734[23] = |(datain[219:216] ^ 0);
  assign w734[24] = |(datain[215:212] ^ 0);
  assign w734[25] = |(datain[211:208] ^ 3);
  assign w734[26] = |(datain[207:204] ^ 14);
  assign w734[27] = |(datain[203:200] ^ 8);
  assign w734[28] = |(datain[199:196] ^ 5);
  assign w734[29] = |(datain[195:192] ^ 14);
  assign w734[30] = |(datain[191:188] ^ 15);
  assign w734[31] = |(datain[187:184] ^ 15);
  assign w734[32] = |(datain[183:180] ^ 12);
  assign w734[33] = |(datain[179:176] ^ 3);
  assign w734[34] = |(datain[175:172] ^ 11);
  assign w734[35] = |(datain[171:168] ^ 4);
  assign w734[36] = |(datain[167:164] ^ 5);
  assign w734[37] = |(datain[163:160] ^ 7);
  assign w734[38] = |(datain[159:156] ^ 2);
  assign w734[39] = |(datain[155:152] ^ 14);
  assign w734[40] = |(datain[151:148] ^ 8);
  assign w734[41] = |(datain[147:144] ^ 11);
  assign w734[42] = |(datain[143:140] ^ 1);
  assign w734[43] = |(datain[139:136] ^ 14);
  assign w734[44] = |(datain[135:132] ^ 15);
  assign w734[45] = |(datain[131:128] ^ 2);
  assign w734[46] = |(datain[127:124] ^ 0);
  assign w734[47] = |(datain[123:120] ^ 2);
  assign w734[48] = |(datain[119:116] ^ 14);
  assign w734[49] = |(datain[115:112] ^ 8);
  assign w734[50] = |(datain[111:108] ^ 5);
  assign w734[51] = |(datain[107:104] ^ 3);
  assign w734[52] = |(datain[103:100] ^ 15);
  assign w734[53] = |(datain[99:96] ^ 15);
  assign w734[54] = |(datain[95:92] ^ 12);
  assign w734[55] = |(datain[91:88] ^ 3);
  assign w734[56] = |(datain[87:84] ^ 11);
  assign w734[57] = |(datain[83:80] ^ 4);
  assign w734[58] = |(datain[79:76] ^ 4);
  assign w734[59] = |(datain[75:72] ^ 0);
  assign w734[60] = |(datain[71:68] ^ 2);
  assign w734[61] = |(datain[67:64] ^ 14);
  assign w734[62] = |(datain[63:60] ^ 8);
  assign w734[63] = |(datain[59:56] ^ 11);
  assign w734[64] = |(datain[55:52] ^ 1);
  assign w734[65] = |(datain[51:48] ^ 14);
  assign w734[66] = |(datain[47:44] ^ 15);
  assign w734[67] = |(datain[43:40] ^ 2);
  assign w734[68] = |(datain[39:36] ^ 0);
  assign w734[69] = |(datain[35:32] ^ 2);
  assign w734[70] = |(datain[31:28] ^ 12);
  assign w734[71] = |(datain[27:24] ^ 13);
  assign w734[72] = |(datain[23:20] ^ 2);
  assign w734[73] = |(datain[19:16] ^ 1);
  assign comp[734] = ~(|w734);
  wire [74-1:0] w735;
  assign w735[0] = |(datain[311:308] ^ 0);
  assign w735[1] = |(datain[307:304] ^ 1);
  assign w735[2] = |(datain[303:300] ^ 11);
  assign w735[3] = |(datain[299:296] ^ 10);
  assign w735[4] = |(datain[295:292] ^ 6);
  assign w735[5] = |(datain[291:288] ^ 9);
  assign w735[6] = |(datain[287:284] ^ 0);
  assign w735[7] = |(datain[283:280] ^ 3);
  assign w735[8] = |(datain[279:276] ^ 12);
  assign w735[9] = |(datain[275:272] ^ 13);
  assign w735[10] = |(datain[271:268] ^ 2);
  assign w735[11] = |(datain[267:264] ^ 1);
  assign w735[12] = |(datain[263:260] ^ 7);
  assign w735[13] = |(datain[259:256] ^ 3);
  assign w735[14] = |(datain[255:252] ^ 0);
  assign w735[15] = |(datain[251:248] ^ 3);
  assign w735[16] = |(datain[247:244] ^ 14);
  assign w735[17] = |(datain[243:240] ^ 9);
  assign w735[18] = |(datain[239:236] ^ 15);
  assign w735[19] = |(datain[235:232] ^ 4);
  assign w735[20] = |(datain[231:228] ^ 15);
  assign w735[21] = |(datain[227:224] ^ 14);
  assign w735[22] = |(datain[223:220] ^ 12);
  assign w735[23] = |(datain[219:216] ^ 3);
  assign w735[24] = |(datain[215:212] ^ 11);
  assign w735[25] = |(datain[211:208] ^ 4);
  assign w735[26] = |(datain[207:204] ^ 5);
  assign w735[27] = |(datain[203:200] ^ 7);
  assign w735[28] = |(datain[199:196] ^ 2);
  assign w735[29] = |(datain[195:192] ^ 14);
  assign w735[30] = |(datain[191:188] ^ 8);
  assign w735[31] = |(datain[187:184] ^ 11);
  assign w735[32] = |(datain[183:180] ^ 1);
  assign w735[33] = |(datain[179:176] ^ 14);
  assign w735[34] = |(datain[175:172] ^ 2);
  assign w735[35] = |(datain[171:168] ^ 15);
  assign w735[36] = |(datain[167:164] ^ 0);
  assign w735[37] = |(datain[163:160] ^ 3);
  assign w735[38] = |(datain[159:156] ^ 12);
  assign w735[39] = |(datain[155:152] ^ 13);
  assign w735[40] = |(datain[151:148] ^ 2);
  assign w735[41] = |(datain[147:144] ^ 1);
  assign w735[42] = |(datain[143:140] ^ 7);
  assign w735[43] = |(datain[139:136] ^ 3);
  assign w735[44] = |(datain[135:132] ^ 0);
  assign w735[45] = |(datain[131:128] ^ 3);
  assign w735[46] = |(datain[127:124] ^ 14);
  assign w735[47] = |(datain[123:120] ^ 9);
  assign w735[48] = |(datain[119:116] ^ 14);
  assign w735[49] = |(datain[115:112] ^ 5);
  assign w735[50] = |(datain[111:108] ^ 15);
  assign w735[51] = |(datain[107:104] ^ 14);
  assign w735[52] = |(datain[103:100] ^ 12);
  assign w735[53] = |(datain[99:96] ^ 3);
  assign w735[54] = |(datain[95:92] ^ 11);
  assign w735[55] = |(datain[91:88] ^ 4);
  assign w735[56] = |(datain[87:84] ^ 4);
  assign w735[57] = |(datain[83:80] ^ 0);
  assign w735[58] = |(datain[79:76] ^ 2);
  assign w735[59] = |(datain[75:72] ^ 14);
  assign w735[60] = |(datain[71:68] ^ 8);
  assign w735[61] = |(datain[67:64] ^ 11);
  assign w735[62] = |(datain[63:60] ^ 1);
  assign w735[63] = |(datain[59:56] ^ 14);
  assign w735[64] = |(datain[55:52] ^ 2);
  assign w735[65] = |(datain[51:48] ^ 15);
  assign w735[66] = |(datain[47:44] ^ 0);
  assign w735[67] = |(datain[43:40] ^ 3);
  assign w735[68] = |(datain[39:36] ^ 12);
  assign w735[69] = |(datain[35:32] ^ 13);
  assign w735[70] = |(datain[31:28] ^ 2);
  assign w735[71] = |(datain[27:24] ^ 1);
  assign w735[72] = |(datain[23:20] ^ 8);
  assign w735[73] = |(datain[19:16] ^ 12);
  assign comp[735] = ~(|w735);
  wire [76-1:0] w736;
  assign w736[0] = |(datain[311:308] ^ 3);
  assign w736[1] = |(datain[307:304] ^ 6);
  assign w736[2] = |(datain[303:300] ^ 3);
  assign w736[3] = |(datain[299:296] ^ 5);
  assign w736[4] = |(datain[295:292] ^ 0);
  assign w736[5] = |(datain[291:288] ^ 4);
  assign w736[6] = |(datain[287:284] ^ 5);
  assign w736[7] = |(datain[283:280] ^ 11);
  assign w736[8] = |(datain[279:276] ^ 12);
  assign w736[9] = |(datain[275:272] ^ 3);
  assign w736[10] = |(datain[271:268] ^ 11);
  assign w736[11] = |(datain[267:264] ^ 9);
  assign w736[12] = |(datain[263:260] ^ 15);
  assign w736[13] = |(datain[259:256] ^ 15);
  assign w736[14] = |(datain[255:252] ^ 0);
  assign w736[15] = |(datain[251:248] ^ 1);
  assign w736[16] = |(datain[247:244] ^ 14);
  assign w736[17] = |(datain[243:240] ^ 8);
  assign w736[18] = |(datain[239:236] ^ 10);
  assign w736[19] = |(datain[235:232] ^ 8);
  assign w736[20] = |(datain[231:228] ^ 15);
  assign w736[21] = |(datain[227:224] ^ 15);
  assign w736[22] = |(datain[223:220] ^ 2);
  assign w736[23] = |(datain[219:216] ^ 14);
  assign w736[24] = |(datain[215:212] ^ 15);
  assign w736[25] = |(datain[211:208] ^ 14);
  assign w736[26] = |(datain[207:204] ^ 0);
  assign w736[27] = |(datain[203:200] ^ 6);
  assign w736[28] = |(datain[199:196] ^ 3);
  assign w736[29] = |(datain[195:192] ^ 5);
  assign w736[30] = |(datain[191:188] ^ 0);
  assign w736[31] = |(datain[187:184] ^ 4);
  assign w736[32] = |(datain[183:180] ^ 14);
  assign w736[33] = |(datain[179:176] ^ 2);
  assign w736[34] = |(datain[175:172] ^ 15);
  assign w736[35] = |(datain[171:168] ^ 6);
  assign w736[36] = |(datain[167:164] ^ 2);
  assign w736[37] = |(datain[163:160] ^ 14);
  assign w736[38] = |(datain[159:156] ^ 15);
  assign w736[39] = |(datain[155:152] ^ 14);
  assign w736[40] = |(datain[151:148] ^ 0);
  assign w736[41] = |(datain[147:144] ^ 14);
  assign w736[42] = |(datain[143:140] ^ 3);
  assign w736[43] = |(datain[139:136] ^ 5);
  assign w736[44] = |(datain[135:132] ^ 0);
  assign w736[45] = |(datain[131:128] ^ 4);
  assign w736[46] = |(datain[127:124] ^ 12);
  assign w736[47] = |(datain[123:120] ^ 3);
  assign w736[48] = |(datain[119:116] ^ 11);
  assign w736[49] = |(datain[115:112] ^ 9);
  assign w736[50] = |(datain[111:108] ^ 15);
  assign w736[51] = |(datain[107:104] ^ 15);
  assign w736[52] = |(datain[103:100] ^ 0);
  assign w736[53] = |(datain[99:96] ^ 1);
  assign w736[54] = |(datain[95:92] ^ 14);
  assign w736[55] = |(datain[91:88] ^ 8);
  assign w736[56] = |(datain[87:84] ^ 9);
  assign w736[57] = |(datain[83:80] ^ 5);
  assign w736[58] = |(datain[79:76] ^ 15);
  assign w736[59] = |(datain[75:72] ^ 15);
  assign w736[60] = |(datain[71:68] ^ 2);
  assign w736[61] = |(datain[67:64] ^ 14);
  assign w736[62] = |(datain[63:60] ^ 15);
  assign w736[63] = |(datain[59:56] ^ 14);
  assign w736[64] = |(datain[55:52] ^ 0);
  assign w736[65] = |(datain[51:48] ^ 14);
  assign w736[66] = |(datain[47:44] ^ 3);
  assign w736[67] = |(datain[43:40] ^ 5);
  assign w736[68] = |(datain[39:36] ^ 0);
  assign w736[69] = |(datain[35:32] ^ 4);
  assign w736[70] = |(datain[31:28] ^ 14);
  assign w736[71] = |(datain[27:24] ^ 2);
  assign w736[72] = |(datain[23:20] ^ 15);
  assign w736[73] = |(datain[19:16] ^ 6);
  assign w736[74] = |(datain[15:12] ^ 12);
  assign w736[75] = |(datain[11:8] ^ 3);
  assign comp[736] = ~(|w736);
  wire [42-1:0] w737;
  assign w737[0] = |(datain[311:308] ^ 11);
  assign w737[1] = |(datain[307:304] ^ 10);
  assign w737[2] = |(datain[303:300] ^ 8);
  assign w737[3] = |(datain[299:296] ^ 5);
  assign w737[4] = |(datain[295:292] ^ 0);
  assign w737[5] = |(datain[291:288] ^ 1);
  assign w737[6] = |(datain[287:284] ^ 11);
  assign w737[7] = |(datain[283:280] ^ 4);
  assign w737[8] = |(datain[279:276] ^ 4);
  assign w737[9] = |(datain[275:272] ^ 14);
  assign w737[10] = |(datain[271:268] ^ 12);
  assign w737[11] = |(datain[267:264] ^ 13);
  assign w737[12] = |(datain[263:260] ^ 2);
  assign w737[13] = |(datain[259:256] ^ 1);
  assign w737[14] = |(datain[255:252] ^ 7);
  assign w737[15] = |(datain[251:248] ^ 2);
  assign w737[16] = |(datain[247:244] ^ 4);
  assign w737[17] = |(datain[243:240] ^ 5);
  assign w737[18] = |(datain[239:236] ^ 11);
  assign w737[19] = |(datain[235:232] ^ 8);
  assign w737[20] = |(datain[231:228] ^ 0);
  assign w737[21] = |(datain[227:224] ^ 0);
  assign w737[22] = |(datain[223:220] ^ 4);
  assign w737[23] = |(datain[219:216] ^ 3);
  assign w737[24] = |(datain[215:212] ^ 11);
  assign w737[25] = |(datain[211:208] ^ 10);
  assign w737[26] = |(datain[207:204] ^ 9);
  assign w737[27] = |(datain[203:200] ^ 14);
  assign w737[28] = |(datain[199:196] ^ 0);
  assign w737[29] = |(datain[195:192] ^ 0);
  assign w737[30] = |(datain[191:188] ^ 12);
  assign w737[31] = |(datain[187:184] ^ 13);
  assign w737[32] = |(datain[183:180] ^ 2);
  assign w737[33] = |(datain[179:176] ^ 1);
  assign w737[34] = |(datain[175:172] ^ 5);
  assign w737[35] = |(datain[171:168] ^ 1);
  assign w737[36] = |(datain[167:164] ^ 11);
  assign w737[37] = |(datain[163:160] ^ 8);
  assign w737[38] = |(datain[159:156] ^ 0);
  assign w737[39] = |(datain[155:152] ^ 1);
  assign w737[40] = |(datain[151:148] ^ 4);
  assign w737[41] = |(datain[147:144] ^ 3);
  assign comp[737] = ~(|w737);
  wire [74-1:0] w738;
  assign w738[0] = |(datain[311:308] ^ 1);
  assign w738[1] = |(datain[307:304] ^ 13);
  assign w738[2] = |(datain[303:300] ^ 8);
  assign w738[3] = |(datain[299:296] ^ 1);
  assign w738[4] = |(datain[295:292] ^ 7);
  assign w738[5] = |(datain[291:288] ^ 15);
  assign w738[6] = |(datain[287:284] ^ 1);
  assign w738[7] = |(datain[283:280] ^ 14);
  assign w738[8] = |(datain[279:276] ^ 4);
  assign w738[9] = |(datain[275:272] ^ 1);
  assign w738[10] = |(datain[271:268] ^ 7);
  assign w738[11] = |(datain[267:264] ^ 4);
  assign w738[12] = |(datain[263:260] ^ 7);
  assign w738[13] = |(datain[259:256] ^ 4);
  assign w738[14] = |(datain[255:252] ^ 1);
  assign w738[15] = |(datain[251:248] ^ 6);
  assign w738[16] = |(datain[247:244] ^ 11);
  assign w738[17] = |(datain[243:240] ^ 1);
  assign w738[18] = |(datain[239:236] ^ 1);
  assign w738[19] = |(datain[235:232] ^ 1);
  assign w738[20] = |(datain[231:228] ^ 8);
  assign w738[21] = |(datain[227:224] ^ 9);
  assign w738[22] = |(datain[223:220] ^ 0);
  assign w738[23] = |(datain[219:216] ^ 14);
  assign w738[24] = |(datain[215:212] ^ 2);
  assign w738[25] = |(datain[211:208] ^ 5);
  assign w738[26] = |(datain[207:204] ^ 0);
  assign w738[27] = |(datain[203:200] ^ 0);
  assign w738[28] = |(datain[199:196] ^ 11);
  assign w738[29] = |(datain[195:192] ^ 8);
  assign w738[30] = |(datain[191:188] ^ 0);
  assign w738[31] = |(datain[187:184] ^ 1);
  assign w738[32] = |(datain[183:180] ^ 0);
  assign w738[33] = |(datain[179:176] ^ 3);
  assign w738[34] = |(datain[175:172] ^ 12);
  assign w738[35] = |(datain[171:168] ^ 13);
  assign w738[36] = |(datain[167:164] ^ 6);
  assign w738[37] = |(datain[163:160] ^ 10);
  assign w738[38] = |(datain[159:156] ^ 7);
  assign w738[39] = |(datain[155:152] ^ 2);
  assign w738[40] = |(datain[151:148] ^ 0);
  assign w738[41] = |(datain[147:144] ^ 9);
  assign w738[42] = |(datain[143:140] ^ 11);
  assign w738[43] = |(datain[139:136] ^ 8);
  assign w738[44] = |(datain[135:132] ^ 0);
  assign w738[45] = |(datain[131:128] ^ 1);
  assign w738[46] = |(datain[127:124] ^ 0);
  assign w738[47] = |(datain[123:120] ^ 3);
  assign w738[48] = |(datain[119:116] ^ 3);
  assign w738[49] = |(datain[115:112] ^ 3);
  assign w738[50] = |(datain[111:108] ^ 13);
  assign w738[51] = |(datain[107:104] ^ 11);
  assign w738[52] = |(datain[103:100] ^ 11);
  assign w738[53] = |(datain[99:96] ^ 1);
  assign w738[54] = |(datain[95:92] ^ 0);
  assign w738[55] = |(datain[91:88] ^ 1);
  assign w738[56] = |(datain[87:84] ^ 12);
  assign w738[57] = |(datain[83:80] ^ 13);
  assign w738[58] = |(datain[79:76] ^ 6);
  assign w738[59] = |(datain[75:72] ^ 10);
  assign w738[60] = |(datain[71:68] ^ 11);
  assign w738[61] = |(datain[67:64] ^ 15);
  assign w738[62] = |(datain[63:60] ^ 3);
  assign w738[63] = |(datain[59:56] ^ 4);
  assign w738[64] = |(datain[55:52] ^ 0);
  assign w738[65] = |(datain[51:48] ^ 0);
  assign w738[66] = |(datain[47:44] ^ 3);
  assign w738[67] = |(datain[43:40] ^ 3);
  assign w738[68] = |(datain[39:36] ^ 13);
  assign w738[69] = |(datain[35:32] ^ 11);
  assign w738[70] = |(datain[31:28] ^ 5);
  assign w738[71] = |(datain[27:24] ^ 3);
  assign w738[72] = |(datain[23:20] ^ 0);
  assign w738[73] = |(datain[19:16] ^ 7);
  assign comp[738] = ~(|w738);
  wire [76-1:0] w739;
  assign w739[0] = |(datain[311:308] ^ 13);
  assign w739[1] = |(datain[307:304] ^ 10);
  assign w739[2] = |(datain[303:300] ^ 9);
  assign w739[3] = |(datain[299:296] ^ 1);
  assign w739[4] = |(datain[295:292] ^ 14);
  assign w739[5] = |(datain[291:288] ^ 8);
  assign w739[6] = |(datain[287:284] ^ 0);
  assign w739[7] = |(datain[283:280] ^ 0);
  assign w739[8] = |(datain[279:276] ^ 0);
  assign w739[9] = |(datain[275:272] ^ 0);
  assign w739[10] = |(datain[271:268] ^ 1);
  assign w739[11] = |(datain[267:264] ^ 0);
  assign w739[12] = |(datain[263:260] ^ 14);
  assign w739[13] = |(datain[259:256] ^ 12);
  assign w739[14] = |(datain[255:252] ^ 3);
  assign w739[15] = |(datain[251:248] ^ 9);
  assign w739[16] = |(datain[247:244] ^ 13);
  assign w739[17] = |(datain[243:240] ^ 0);
  assign w739[18] = |(datain[239:236] ^ 14);
  assign w739[19] = |(datain[235:232] ^ 10);
  assign w739[20] = |(datain[231:228] ^ 11);
  assign w739[21] = |(datain[227:224] ^ 4);
  assign w739[22] = |(datain[223:220] ^ 3);
  assign w739[23] = |(datain[219:216] ^ 3);
  assign w739[24] = |(datain[215:212] ^ 0);
  assign w739[25] = |(datain[211:208] ^ 0);
  assign w739[26] = |(datain[207:204] ^ 3);
  assign w739[27] = |(datain[203:200] ^ 0);
  assign w739[28] = |(datain[199:196] ^ 14);
  assign w739[29] = |(datain[195:192] ^ 10);
  assign w739[30] = |(datain[191:188] ^ 6);
  assign w739[31] = |(datain[187:184] ^ 6);
  assign w739[32] = |(datain[183:180] ^ 7);
  assign w739[33] = |(datain[179:176] ^ 6);
  assign w739[34] = |(datain[175:172] ^ 10);
  assign w739[35] = |(datain[171:168] ^ 4);
  assign w739[36] = |(datain[167:164] ^ 14);
  assign w739[37] = |(datain[163:160] ^ 8);
  assign w739[38] = |(datain[159:156] ^ 0);
  assign w739[39] = |(datain[155:152] ^ 0);
  assign w739[40] = |(datain[151:148] ^ 0);
  assign w739[41] = |(datain[147:144] ^ 0);
  assign w739[42] = |(datain[143:140] ^ 1);
  assign w739[43] = |(datain[139:136] ^ 0);
  assign w739[44] = |(datain[135:132] ^ 14);
  assign w739[45] = |(datain[131:128] ^ 11);
  assign w739[46] = |(datain[127:124] ^ 6);
  assign w739[47] = |(datain[123:120] ^ 3);
  assign w739[48] = |(datain[119:116] ^ 9);
  assign w739[49] = |(datain[115:112] ^ 6);
  assign w739[50] = |(datain[111:108] ^ 15);
  assign w739[51] = |(datain[107:104] ^ 5);
  assign w739[52] = |(datain[103:100] ^ 11);
  assign w739[53] = |(datain[99:96] ^ 9);
  assign w739[54] = |(datain[95:92] ^ 5);
  assign w739[55] = |(datain[91:88] ^ 5);
  assign w739[56] = |(datain[87:84] ^ 0);
  assign w739[57] = |(datain[83:80] ^ 0);
  assign w739[58] = |(datain[79:76] ^ 3);
  assign w739[59] = |(datain[75:72] ^ 0);
  assign w739[60] = |(datain[71:68] ^ 4);
  assign w739[61] = |(datain[67:64] ^ 7);
  assign w739[62] = |(datain[63:60] ^ 13);
  assign w739[63] = |(datain[59:56] ^ 10);
  assign w739[64] = |(datain[55:52] ^ 7);
  assign w739[65] = |(datain[51:48] ^ 1);
  assign w739[66] = |(datain[47:44] ^ 1);
  assign w739[67] = |(datain[43:40] ^ 5);
  assign w739[68] = |(datain[39:36] ^ 14);
  assign w739[69] = |(datain[35:32] ^ 8);
  assign w739[70] = |(datain[31:28] ^ 0);
  assign w739[71] = |(datain[27:24] ^ 0);
  assign w739[72] = |(datain[23:20] ^ 0);
  assign w739[73] = |(datain[19:16] ^ 0);
  assign w739[74] = |(datain[15:12] ^ 1);
  assign w739[75] = |(datain[11:8] ^ 0);
  assign comp[739] = ~(|w739);
  wire [54-1:0] w740;
  assign w740[0] = |(datain[311:308] ^ 5);
  assign w740[1] = |(datain[307:304] ^ 13);
  assign w740[2] = |(datain[303:300] ^ 8);
  assign w740[3] = |(datain[299:296] ^ 1);
  assign w740[4] = |(datain[295:292] ^ 14);
  assign w740[5] = |(datain[291:288] ^ 13);
  assign w740[6] = |(datain[287:284] ^ 0);
  assign w740[7] = |(datain[283:280] ^ 10);
  assign w740[8] = |(datain[279:276] ^ 0);
  assign w740[9] = |(datain[275:272] ^ 1);
  assign w740[10] = |(datain[271:268] ^ 8);
  assign w740[11] = |(datain[267:264] ^ 13);
  assign w740[12] = |(datain[263:260] ^ 11);
  assign w740[13] = |(datain[259:256] ^ 6);
  assign w740[14] = |(datain[255:252] ^ 2);
  assign w740[15] = |(datain[251:248] ^ 5);
  assign w740[16] = |(datain[247:244] ^ 0);
  assign w740[17] = |(datain[243:240] ^ 1);
  assign w740[18] = |(datain[239:236] ^ 5);
  assign w740[19] = |(datain[235:232] ^ 6);
  assign w740[20] = |(datain[231:228] ^ 8);
  assign w740[21] = |(datain[227:224] ^ 11);
  assign w740[22] = |(datain[223:220] ^ 15);
  assign w740[23] = |(datain[219:216] ^ 14);
  assign w740[24] = |(datain[215:212] ^ 8);
  assign w740[25] = |(datain[211:208] ^ 11);
  assign w740[26] = |(datain[207:204] ^ 9);
  assign w740[27] = |(datain[203:200] ^ 6);
  assign w740[28] = |(datain[199:196] ^ 8);
  assign w740[29] = |(datain[195:192] ^ 13);
  assign w740[30] = |(datain[191:188] ^ 0);
  assign w740[31] = |(datain[187:184] ^ 2);
  assign w740[32] = |(datain[183:180] ^ 11);
  assign w740[33] = |(datain[179:176] ^ 9);
  assign w740[34] = |(datain[175:172] ^ 6);
  assign w740[35] = |(datain[171:168] ^ 8);
  assign w740[36] = |(datain[167:164] ^ 0);
  assign w740[37] = |(datain[163:160] ^ 1);
  assign w740[38] = |(datain[159:156] ^ 15);
  assign w740[39] = |(datain[155:152] ^ 12);
  assign w740[40] = |(datain[151:148] ^ 10);
  assign w740[41] = |(datain[147:144] ^ 12);
  assign w740[42] = |(datain[143:140] ^ 3);
  assign w740[43] = |(datain[139:136] ^ 2);
  assign w740[44] = |(datain[135:132] ^ 12);
  assign w740[45] = |(datain[131:128] ^ 2);
  assign w740[46] = |(datain[127:124] ^ 10);
  assign w740[47] = |(datain[123:120] ^ 10);
  assign w740[48] = |(datain[119:116] ^ 14);
  assign w740[49] = |(datain[115:112] ^ 2);
  assign w740[50] = |(datain[111:108] ^ 15);
  assign w740[51] = |(datain[107:104] ^ 10);
  assign w740[52] = |(datain[103:100] ^ 12);
  assign w740[53] = |(datain[99:96] ^ 3);
  assign comp[740] = ~(|w740);
  wire [42-1:0] w741;
  assign w741[0] = |(datain[311:308] ^ 0);
  assign w741[1] = |(datain[307:304] ^ 2);
  assign w741[2] = |(datain[303:300] ^ 8);
  assign w741[3] = |(datain[299:296] ^ 11);
  assign w741[4] = |(datain[295:292] ^ 15);
  assign w741[5] = |(datain[291:288] ^ 2);
  assign w741[6] = |(datain[287:284] ^ 8);
  assign w741[7] = |(datain[283:280] ^ 10);
  assign w741[8] = |(datain[279:276] ^ 2);
  assign w741[9] = |(datain[275:272] ^ 3);
  assign w741[10] = |(datain[271:268] ^ 8);
  assign w741[11] = |(datain[267:264] ^ 11);
  assign w741[12] = |(datain[263:260] ^ 1);
  assign w741[13] = |(datain[259:256] ^ 6);
  assign w741[14] = |(datain[255:252] ^ 3);
  assign w741[15] = |(datain[251:248] ^ 14);
  assign w741[16] = |(datain[247:244] ^ 0);
  assign w741[17] = |(datain[243:240] ^ 15);
  assign w741[18] = |(datain[239:236] ^ 15);
  assign w741[19] = |(datain[235:232] ^ 12);
  assign w741[20] = |(datain[231:228] ^ 14);
  assign w741[21] = |(datain[227:224] ^ 11);
  assign w741[22] = |(datain[223:220] ^ 4);
  assign w741[23] = |(datain[219:216] ^ 5);
  assign w741[24] = |(datain[215:212] ^ 9);
  assign w741[25] = |(datain[211:208] ^ 0);
  assign w741[26] = |(datain[207:204] ^ 12);
  assign w741[27] = |(datain[203:200] ^ 13);
  assign w741[28] = |(datain[199:196] ^ 1);
  assign w741[29] = |(datain[195:192] ^ 3);
  assign w741[30] = |(datain[191:188] ^ 8);
  assign w741[31] = |(datain[187:184] ^ 10);
  assign w741[32] = |(datain[183:180] ^ 2);
  assign w741[33] = |(datain[179:176] ^ 2);
  assign w741[34] = |(datain[175:172] ^ 11);
  assign w741[35] = |(datain[171:168] ^ 4);
  assign w741[36] = |(datain[167:164] ^ 0);
  assign w741[37] = |(datain[163:160] ^ 0);
  assign w741[38] = |(datain[159:156] ^ 8);
  assign w741[39] = |(datain[155:152] ^ 1);
  assign w741[40] = |(datain[151:148] ^ 14);
  assign w741[41] = |(datain[147:144] ^ 1);
  assign comp[741] = ~(|w741);
  wire [32-1:0] w742;
  assign w742[0] = |(datain[311:308] ^ 0);
  assign w742[1] = |(datain[307:304] ^ 1);
  assign w742[2] = |(datain[303:300] ^ 9);
  assign w742[3] = |(datain[299:296] ^ 0);
  assign w742[4] = |(datain[295:292] ^ 14);
  assign w742[5] = |(datain[291:288] ^ 8);
  assign w742[6] = |(datain[287:284] ^ 0);
  assign w742[7] = |(datain[283:280] ^ 0);
  assign w742[8] = |(datain[279:276] ^ 0);
  assign w742[9] = |(datain[275:272] ^ 0);
  assign w742[10] = |(datain[271:268] ^ 5);
  assign w742[11] = |(datain[267:264] ^ 14);
  assign w742[12] = |(datain[263:260] ^ 5);
  assign w742[13] = |(datain[259:256] ^ 6);
  assign w742[14] = |(datain[255:252] ^ 11);
  assign w742[15] = |(datain[251:248] ^ 10);
  assign w742[16] = |(datain[247:244] ^ 4);
  assign w742[17] = |(datain[243:240] ^ 12);
  assign w742[18] = |(datain[239:236] ^ 0);
  assign w742[19] = |(datain[235:232] ^ 8);
  assign w742[20] = |(datain[231:228] ^ 8);
  assign w742[21] = |(datain[227:224] ^ 1);
  assign w742[22] = |(datain[223:220] ^ 14);
  assign w742[23] = |(datain[219:216] ^ 10);
  assign w742[24] = |(datain[215:212] ^ 0);
  assign w742[25] = |(datain[211:208] ^ 0);
  assign w742[26] = |(datain[207:204] ^ 0);
  assign w742[27] = |(datain[203:200] ^ 1);
  assign w742[28] = |(datain[199:196] ^ 8);
  assign w742[29] = |(datain[195:192] ^ 3);
  assign w742[30] = |(datain[191:188] ^ 14);
  assign w742[31] = |(datain[187:184] ^ 14);
  assign comp[742] = ~(|w742);
  wire [28-1:0] w743;
  assign w743[0] = |(datain[311:308] ^ 9);
  assign w743[1] = |(datain[307:304] ^ 0);
  assign w743[2] = |(datain[303:300] ^ 14);
  assign w743[3] = |(datain[299:296] ^ 8);
  assign w743[4] = |(datain[295:292] ^ 0);
  assign w743[5] = |(datain[291:288] ^ 0);
  assign w743[6] = |(datain[287:284] ^ 0);
  assign w743[7] = |(datain[283:280] ^ 0);
  assign w743[8] = |(datain[279:276] ^ 5);
  assign w743[9] = |(datain[275:272] ^ 14);
  assign w743[10] = |(datain[271:268] ^ 5);
  assign w743[11] = |(datain[267:264] ^ 6);
  assign w743[12] = |(datain[263:260] ^ 11);
  assign w743[13] = |(datain[259:256] ^ 10);
  assign w743[14] = |(datain[255:252] ^ 4);
  assign w743[15] = |(datain[251:248] ^ 12);
  assign w743[16] = |(datain[247:244] ^ 0);
  assign w743[17] = |(datain[243:240] ^ 8);
  assign w743[18] = |(datain[239:236] ^ 8);
  assign w743[19] = |(datain[235:232] ^ 1);
  assign w743[20] = |(datain[231:228] ^ 14);
  assign w743[21] = |(datain[227:224] ^ 10);
  assign w743[22] = |(datain[223:220] ^ 0);
  assign w743[23] = |(datain[219:216] ^ 0);
  assign w743[24] = |(datain[215:212] ^ 0);
  assign w743[25] = |(datain[211:208] ^ 1);
  assign w743[26] = |(datain[207:204] ^ 8);
  assign w743[27] = |(datain[203:200] ^ 3);
  assign comp[743] = ~(|w743);
  wire [60-1:0] w744;
  assign w744[0] = |(datain[311:308] ^ 14);
  assign w744[1] = |(datain[307:304] ^ 8);
  assign w744[2] = |(datain[303:300] ^ 0);
  assign w744[3] = |(datain[299:296] ^ 0);
  assign w744[4] = |(datain[295:292] ^ 0);
  assign w744[5] = |(datain[291:288] ^ 0);
  assign w744[6] = |(datain[287:284] ^ 5);
  assign w744[7] = |(datain[283:280] ^ 13);
  assign w744[8] = |(datain[279:276] ^ 8);
  assign w744[9] = |(datain[275:272] ^ 1);
  assign w744[10] = |(datain[271:268] ^ 14);
  assign w744[11] = |(datain[267:264] ^ 13);
  assign w744[12] = |(datain[263:260] ^ 0);
  assign w744[13] = |(datain[259:256] ^ 10);
  assign w744[14] = |(datain[255:252] ^ 0);
  assign w744[15] = |(datain[251:248] ^ 1);
  assign w744[16] = |(datain[247:244] ^ 8);
  assign w744[17] = |(datain[243:240] ^ 13);
  assign w744[18] = |(datain[239:236] ^ 11);
  assign w744[19] = |(datain[235:232] ^ 6);
  assign w744[20] = |(datain[231:228] ^ 2);
  assign w744[21] = |(datain[227:224] ^ 5);
  assign w744[22] = |(datain[223:220] ^ 0);
  assign w744[23] = |(datain[219:216] ^ 1);
  assign w744[24] = |(datain[215:212] ^ 5);
  assign w744[25] = |(datain[211:208] ^ 6);
  assign w744[26] = |(datain[207:204] ^ 8);
  assign w744[27] = |(datain[203:200] ^ 11);
  assign w744[28] = |(datain[199:196] ^ 15);
  assign w744[29] = |(datain[195:192] ^ 14);
  assign w744[30] = |(datain[191:188] ^ 8);
  assign w744[31] = |(datain[187:184] ^ 11);
  assign w744[32] = |(datain[183:180] ^ 9);
  assign w744[33] = |(datain[179:176] ^ 6);
  assign w744[34] = |(datain[175:172] ^ 8);
  assign w744[35] = |(datain[171:168] ^ 3);
  assign w744[36] = |(datain[167:164] ^ 0);
  assign w744[37] = |(datain[163:160] ^ 2);
  assign w744[38] = |(datain[159:156] ^ 11);
  assign w744[39] = |(datain[155:152] ^ 9);
  assign w744[40] = |(datain[151:148] ^ 5);
  assign w744[41] = |(datain[147:144] ^ 14);
  assign w744[42] = |(datain[143:140] ^ 0);
  assign w744[43] = |(datain[139:136] ^ 1);
  assign w744[44] = |(datain[135:132] ^ 15);
  assign w744[45] = |(datain[131:128] ^ 12);
  assign w744[46] = |(datain[127:124] ^ 10);
  assign w744[47] = |(datain[123:120] ^ 12);
  assign w744[48] = |(datain[119:116] ^ 3);
  assign w744[49] = |(datain[115:112] ^ 2);
  assign w744[50] = |(datain[111:108] ^ 12);
  assign w744[51] = |(datain[107:104] ^ 2);
  assign w744[52] = |(datain[103:100] ^ 10);
  assign w744[53] = |(datain[99:96] ^ 10);
  assign w744[54] = |(datain[95:92] ^ 14);
  assign w744[55] = |(datain[91:88] ^ 2);
  assign w744[56] = |(datain[87:84] ^ 15);
  assign w744[57] = |(datain[83:80] ^ 10);
  assign w744[58] = |(datain[79:76] ^ 12);
  assign w744[59] = |(datain[75:72] ^ 3);
  assign comp[744] = ~(|w744);
  wire [46-1:0] w745;
  assign w745[0] = |(datain[311:308] ^ 12);
  assign w745[1] = |(datain[307:304] ^ 0);
  assign w745[2] = |(datain[303:300] ^ 8);
  assign w745[3] = |(datain[299:296] ^ 14);
  assign w745[4] = |(datain[295:292] ^ 13);
  assign w745[5] = |(datain[291:288] ^ 8);
  assign w745[6] = |(datain[287:284] ^ 8);
  assign w745[7] = |(datain[283:280] ^ 1);
  assign w745[8] = |(datain[279:276] ^ 3);
  assign w745[9] = |(datain[275:272] ^ 15);
  assign w745[10] = |(datain[271:268] ^ 15);
  assign w745[11] = |(datain[267:264] ^ 15);
  assign w745[12] = |(datain[263:260] ^ 1);
  assign w745[13] = |(datain[259:256] ^ 0);
  assign w745[14] = |(datain[255:252] ^ 7);
  assign w745[15] = |(datain[251:248] ^ 4);
  assign w745[16] = |(datain[247:244] ^ 2);
  assign w745[17] = |(datain[243:240] ^ 5);
  assign w745[18] = |(datain[239:236] ^ 12);
  assign w745[19] = |(datain[235:232] ^ 7);
  assign w745[20] = |(datain[231:228] ^ 0);
  assign w745[21] = |(datain[227:224] ^ 7);
  assign w745[22] = |(datain[223:220] ^ 15);
  assign w745[23] = |(datain[219:216] ^ 15);
  assign w745[24] = |(datain[215:212] ^ 1);
  assign w745[25] = |(datain[211:208] ^ 0);
  assign w745[26] = |(datain[207:204] ^ 1);
  assign w745[27] = |(datain[203:200] ^ 15);
  assign w745[28] = |(datain[199:196] ^ 15);
  assign w745[29] = |(datain[195:192] ^ 12);
  assign w745[30] = |(datain[191:188] ^ 15);
  assign w745[31] = |(datain[187:184] ^ 3);
  assign w745[32] = |(datain[183:180] ^ 10);
  assign w745[33] = |(datain[179:176] ^ 4);
  assign w745[34] = |(datain[175:172] ^ 2);
  assign w745[35] = |(datain[171:168] ^ 14);
  assign w745[36] = |(datain[167:164] ^ 8);
  assign w745[37] = |(datain[163:160] ^ 11);
  assign w745[38] = |(datain[159:156] ^ 1);
  assign w745[39] = |(datain[155:152] ^ 14);
  assign w745[40] = |(datain[151:148] ^ 13);
  assign w745[41] = |(datain[147:144] ^ 5);
  assign w745[42] = |(datain[143:140] ^ 0);
  assign w745[43] = |(datain[139:136] ^ 2);
  assign w745[44] = |(datain[135:132] ^ 8);
  assign w745[45] = |(datain[131:128] ^ 14);
  assign comp[745] = ~(|w745);
  wire [46-1:0] w746;
  assign w746[0] = |(datain[311:308] ^ 6);
  assign w746[1] = |(datain[307:304] ^ 3);
  assign w746[2] = |(datain[303:300] ^ 0);
  assign w746[3] = |(datain[299:296] ^ 6);
  assign w746[4] = |(datain[295:292] ^ 8);
  assign w746[5] = |(datain[291:288] ^ 12);
  assign w746[6] = |(datain[287:284] ^ 12);
  assign w746[7] = |(datain[283:280] ^ 8);
  assign w746[8] = |(datain[279:276] ^ 8);
  assign w746[9] = |(datain[275:272] ^ 14);
  assign w746[10] = |(datain[271:268] ^ 13);
  assign w746[11] = |(datain[267:264] ^ 8);
  assign w746[12] = |(datain[263:260] ^ 11);
  assign w746[13] = |(datain[259:256] ^ 15);
  assign w746[14] = |(datain[255:252] ^ 0);
  assign w746[15] = |(datain[251:248] ^ 0);
  assign w746[16] = |(datain[247:244] ^ 0);
  assign w746[17] = |(datain[243:240] ^ 0);
  assign w746[18] = |(datain[239:236] ^ 11);
  assign w746[19] = |(datain[235:232] ^ 8);
  assign w746[20] = |(datain[231:228] ^ 6);
  assign w746[21] = |(datain[227:224] ^ 0);
  assign w746[22] = |(datain[223:220] ^ 9);
  assign w746[23] = |(datain[219:216] ^ 15);
  assign w746[24] = |(datain[215:212] ^ 8);
  assign w746[25] = |(datain[211:208] ^ 14);
  assign w746[26] = |(datain[207:204] ^ 12);
  assign w746[27] = |(datain[203:200] ^ 0);
  assign w746[28] = |(datain[199:196] ^ 11);
  assign w746[29] = |(datain[195:192] ^ 14);
  assign w746[30] = |(datain[191:188] ^ 0);
  assign w746[31] = |(datain[187:184] ^ 0);
  assign w746[32] = |(datain[183:180] ^ 0);
  assign w746[33] = |(datain[179:176] ^ 0);
  assign w746[34] = |(datain[175:172] ^ 11);
  assign w746[35] = |(datain[171:168] ^ 11);
  assign w746[36] = |(datain[167:164] ^ 0);
  assign w746[37] = |(datain[163:160] ^ 7);
  assign w746[38] = |(datain[159:156] ^ 0);
  assign w746[39] = |(datain[155:152] ^ 2);
  assign w746[40] = |(datain[151:148] ^ 2);
  assign w746[41] = |(datain[147:144] ^ 6);
  assign w746[42] = |(datain[143:140] ^ 8);
  assign w746[43] = |(datain[139:136] ^ 11);
  assign w746[44] = |(datain[135:132] ^ 0);
  assign w746[45] = |(datain[131:128] ^ 7);
  assign comp[746] = ~(|w746);
  wire [48-1:0] w747;
  assign w747[0] = |(datain[311:308] ^ 5);
  assign w747[1] = |(datain[307:304] ^ 6);
  assign w747[2] = |(datain[303:300] ^ 1);
  assign w747[3] = |(datain[299:296] ^ 13);
  assign w747[4] = |(datain[295:292] ^ 12);
  assign w747[5] = |(datain[291:288] ^ 7);
  assign w747[6] = |(datain[287:284] ^ 12);
  assign w747[7] = |(datain[283:280] ^ 4);
  assign w747[8] = |(datain[279:276] ^ 1);
  assign w747[9] = |(datain[275:272] ^ 0);
  assign w747[10] = |(datain[271:268] ^ 7);
  assign w747[11] = |(datain[267:264] ^ 11);
  assign w747[12] = |(datain[263:260] ^ 5);
  assign w747[13] = |(datain[259:256] ^ 5);
  assign w747[14] = |(datain[255:252] ^ 2);
  assign w747[15] = |(datain[251:248] ^ 7);
  assign w747[16] = |(datain[247:244] ^ 12);
  assign w747[17] = |(datain[243:240] ^ 3);
  assign w747[18] = |(datain[239:236] ^ 8);
  assign w747[19] = |(datain[235:232] ^ 12);
  assign w747[20] = |(datain[231:228] ^ 8);
  assign w747[21] = |(datain[227:224] ^ 12);
  assign w747[22] = |(datain[223:220] ^ 14);
  assign w747[23] = |(datain[219:216] ^ 3);
  assign w747[24] = |(datain[215:212] ^ 0);
  assign w747[25] = |(datain[211:208] ^ 0);
  assign w747[26] = |(datain[207:204] ^ 10);
  assign w747[27] = |(datain[203:200] ^ 2);
  assign w747[28] = |(datain[199:196] ^ 14);
  assign w747[29] = |(datain[195:192] ^ 2);
  assign w747[30] = |(datain[191:188] ^ 11);
  assign w747[31] = |(datain[187:184] ^ 6);
  assign w747[32] = |(datain[183:180] ^ 2);
  assign w747[33] = |(datain[179:176] ^ 14);
  assign w747[34] = |(datain[175:172] ^ 14);
  assign w747[35] = |(datain[171:168] ^ 8);
  assign w747[36] = |(datain[167:164] ^ 6);
  assign w747[37] = |(datain[163:160] ^ 15);
  assign w747[38] = |(datain[159:156] ^ 6);
  assign w747[39] = |(datain[155:152] ^ 8);
  assign w747[40] = |(datain[151:148] ^ 10);
  assign w747[41] = |(datain[147:144] ^ 8);
  assign w747[42] = |(datain[143:140] ^ 11);
  assign w747[43] = |(datain[139:136] ^ 15);
  assign w747[44] = |(datain[135:132] ^ 9);
  assign w747[45] = |(datain[131:128] ^ 8);
  assign w747[46] = |(datain[127:124] ^ 1);
  assign w747[47] = |(datain[123:120] ^ 10);
  assign comp[747] = ~(|w747);
  wire [48-1:0] w748;
  assign w748[0] = |(datain[311:308] ^ 2);
  assign w748[1] = |(datain[307:304] ^ 0);
  assign w748[2] = |(datain[303:300] ^ 13);
  assign w748[3] = |(datain[299:296] ^ 2);
  assign w748[4] = |(datain[295:292] ^ 7);
  assign w748[5] = |(datain[291:288] ^ 4);
  assign w748[6] = |(datain[287:284] ^ 8);
  assign w748[7] = |(datain[283:280] ^ 8);
  assign w748[8] = |(datain[279:276] ^ 7);
  assign w748[9] = |(datain[275:272] ^ 11);
  assign w748[10] = |(datain[271:268] ^ 14);
  assign w748[11] = |(datain[267:264] ^ 6);
  assign w748[12] = |(datain[263:260] ^ 9);
  assign w748[13] = |(datain[259:256] ^ 12);
  assign w748[14] = |(datain[255:252] ^ 15);
  assign w748[15] = |(datain[251:248] ^ 2);
  assign w748[16] = |(datain[247:244] ^ 7);
  assign w748[17] = |(datain[243:240] ^ 1);
  assign w748[18] = |(datain[239:236] ^ 10);
  assign w748[19] = |(datain[235:232] ^ 15);
  assign w748[20] = |(datain[231:228] ^ 6);
  assign w748[21] = |(datain[227:224] ^ 2);
  assign w748[22] = |(datain[223:220] ^ 1);
  assign w748[23] = |(datain[219:216] ^ 3);
  assign w748[24] = |(datain[215:212] ^ 15);
  assign w748[25] = |(datain[211:208] ^ 13);
  assign w748[26] = |(datain[207:204] ^ 3);
  assign w748[27] = |(datain[203:200] ^ 8);
  assign w748[28] = |(datain[199:196] ^ 11);
  assign w748[29] = |(datain[195:192] ^ 1);
  assign w748[30] = |(datain[191:188] ^ 6);
  assign w748[31] = |(datain[187:184] ^ 9);
  assign w748[32] = |(datain[183:180] ^ 6);
  assign w748[33] = |(datain[179:176] ^ 0);
  assign w748[34] = |(datain[175:172] ^ 13);
  assign w748[35] = |(datain[171:168] ^ 7);
  assign w748[36] = |(datain[167:164] ^ 4);
  assign w748[37] = |(datain[163:160] ^ 12);
  assign w748[38] = |(datain[159:156] ^ 10);
  assign w748[39] = |(datain[155:152] ^ 4);
  assign w748[40] = |(datain[151:148] ^ 7);
  assign w748[41] = |(datain[147:144] ^ 11);
  assign w748[42] = |(datain[143:140] ^ 1);
  assign w748[43] = |(datain[139:136] ^ 14);
  assign w748[44] = |(datain[135:132] ^ 6);
  assign w748[45] = |(datain[131:128] ^ 15);
  assign w748[46] = |(datain[127:124] ^ 6);
  assign w748[47] = |(datain[123:120] ^ 14);
  assign comp[748] = ~(|w748);
  wire [74-1:0] w749;
  assign w749[0] = |(datain[311:308] ^ 1);
  assign w749[1] = |(datain[307:304] ^ 12);
  assign w749[2] = |(datain[303:300] ^ 0);
  assign w749[3] = |(datain[299:296] ^ 0);
  assign w749[4] = |(datain[295:292] ^ 8);
  assign w749[5] = |(datain[291:288] ^ 13);
  assign w749[6] = |(datain[287:284] ^ 1);
  assign w749[7] = |(datain[283:280] ^ 6);
  assign w749[8] = |(datain[279:276] ^ 0);
  assign w749[9] = |(datain[275:272] ^ 3);
  assign w749[10] = |(datain[271:268] ^ 0);
  assign w749[11] = |(datain[267:264] ^ 1);
  assign w749[12] = |(datain[263:260] ^ 11);
  assign w749[13] = |(datain[259:256] ^ 4);
  assign w749[14] = |(datain[255:252] ^ 4);
  assign w749[15] = |(datain[251:248] ^ 0);
  assign w749[16] = |(datain[247:244] ^ 12);
  assign w749[17] = |(datain[243:240] ^ 13);
  assign w749[18] = |(datain[239:236] ^ 2);
  assign w749[19] = |(datain[235:232] ^ 1);
  assign w749[20] = |(datain[231:228] ^ 7);
  assign w749[21] = |(datain[227:224] ^ 2);
  assign w749[22] = |(datain[223:220] ^ 1);
  assign w749[23] = |(datain[219:216] ^ 0);
  assign w749[24] = |(datain[215:212] ^ 14);
  assign w749[25] = |(datain[211:208] ^ 8);
  assign w749[26] = |(datain[207:204] ^ 7);
  assign w749[27] = |(datain[203:200] ^ 13);
  assign w749[28] = |(datain[199:196] ^ 0);
  assign w749[29] = |(datain[195:192] ^ 0);
  assign w749[30] = |(datain[191:188] ^ 7);
  assign w749[31] = |(datain[187:184] ^ 2);
  assign w749[32] = |(datain[183:180] ^ 0);
  assign w749[33] = |(datain[179:176] ^ 11);
  assign w749[34] = |(datain[175:172] ^ 11);
  assign w749[35] = |(datain[171:168] ^ 9);
  assign w749[36] = |(datain[167:164] ^ 6);
  assign w749[37] = |(datain[163:160] ^ 7);
  assign w749[38] = |(datain[159:156] ^ 0);
  assign w749[39] = |(datain[155:152] ^ 4);
  assign w749[40] = |(datain[151:148] ^ 8);
  assign w749[41] = |(datain[147:144] ^ 13);
  assign w749[42] = |(datain[143:140] ^ 1);
  assign w749[43] = |(datain[139:136] ^ 6);
  assign w749[44] = |(datain[135:132] ^ 0);
  assign w749[45] = |(datain[131:128] ^ 0);
  assign w749[46] = |(datain[127:124] ^ 0);
  assign w749[47] = |(datain[123:120] ^ 1);
  assign w749[48] = |(datain[119:116] ^ 11);
  assign w749[49] = |(datain[115:112] ^ 4);
  assign w749[50] = |(datain[111:108] ^ 4);
  assign w749[51] = |(datain[107:104] ^ 0);
  assign w749[52] = |(datain[103:100] ^ 12);
  assign w749[53] = |(datain[99:96] ^ 13);
  assign w749[54] = |(datain[95:92] ^ 2);
  assign w749[55] = |(datain[91:88] ^ 1);
  assign w749[56] = |(datain[87:84] ^ 2);
  assign w749[57] = |(datain[83:80] ^ 14);
  assign w749[58] = |(datain[79:76] ^ 8);
  assign w749[59] = |(datain[75:72] ^ 11);
  assign w749[60] = |(datain[71:68] ^ 1);
  assign w749[61] = |(datain[67:64] ^ 14);
  assign w749[62] = |(datain[63:60] ^ 5);
  assign w749[63] = |(datain[59:56] ^ 4);
  assign w749[64] = |(datain[55:52] ^ 0);
  assign w749[65] = |(datain[51:48] ^ 1);
  assign w749[66] = |(datain[47:44] ^ 2);
  assign w749[67] = |(datain[43:40] ^ 14);
  assign w749[68] = |(datain[39:36] ^ 8);
  assign w749[69] = |(datain[35:32] ^ 11);
  assign w749[70] = |(datain[31:28] ^ 1);
  assign w749[71] = |(datain[27:24] ^ 6);
  assign w749[72] = |(datain[23:20] ^ 4);
  assign w749[73] = |(datain[19:16] ^ 12);
  assign comp[749] = ~(|w749);
  wire [74-1:0] w750;
  assign w750[0] = |(datain[311:308] ^ 0);
  assign w750[1] = |(datain[307:304] ^ 1);
  assign w750[2] = |(datain[303:300] ^ 7);
  assign w750[3] = |(datain[299:296] ^ 3);
  assign w750[4] = |(datain[295:292] ^ 0);
  assign w750[5] = |(datain[291:288] ^ 3);
  assign w750[6] = |(datain[287:284] ^ 14);
  assign w750[7] = |(datain[283:280] ^ 9);
  assign w750[8] = |(datain[279:276] ^ 15);
  assign w750[9] = |(datain[275:272] ^ 13);
  assign w750[10] = |(datain[271:268] ^ 0);
  assign w750[11] = |(datain[267:264] ^ 0);
  assign w750[12] = |(datain[263:260] ^ 11);
  assign w750[13] = |(datain[259:256] ^ 9);
  assign w750[14] = |(datain[255:252] ^ 0);
  assign w750[15] = |(datain[251:248] ^ 3);
  assign w750[16] = |(datain[247:244] ^ 0);
  assign w750[17] = |(datain[243:240] ^ 0);
  assign w750[18] = |(datain[239:236] ^ 8);
  assign w750[19] = |(datain[235:232] ^ 13);
  assign w750[20] = |(datain[231:228] ^ 1);
  assign w750[21] = |(datain[227:224] ^ 6);
  assign w750[22] = |(datain[223:220] ^ 2);
  assign w750[23] = |(datain[219:216] ^ 4);
  assign w750[24] = |(datain[215:212] ^ 0);
  assign w750[25] = |(datain[211:208] ^ 1);
  assign w750[26] = |(datain[207:204] ^ 11);
  assign w750[27] = |(datain[203:200] ^ 4);
  assign w750[28] = |(datain[199:196] ^ 4);
  assign w750[29] = |(datain[195:192] ^ 0);
  assign w750[30] = |(datain[191:188] ^ 12);
  assign w750[31] = |(datain[187:184] ^ 13);
  assign w750[32] = |(datain[183:180] ^ 2);
  assign w750[33] = |(datain[179:176] ^ 1);
  assign w750[34] = |(datain[175:172] ^ 14);
  assign w750[35] = |(datain[171:168] ^ 9);
  assign w750[36] = |(datain[167:164] ^ 14);
  assign w750[37] = |(datain[163:160] ^ 15);
  assign w750[38] = |(datain[159:156] ^ 0);
  assign w750[39] = |(datain[155:152] ^ 0);
  assign w750[40] = |(datain[151:148] ^ 0);
  assign w750[41] = |(datain[147:144] ^ 14);
  assign w750[42] = |(datain[143:140] ^ 1);
  assign w750[43] = |(datain[139:136] ^ 15);
  assign w750[44] = |(datain[135:132] ^ 14);
  assign w750[45] = |(datain[131:128] ^ 8);
  assign w750[46] = |(datain[127:124] ^ 4);
  assign w750[47] = |(datain[123:120] ^ 11);
  assign w750[48] = |(datain[119:116] ^ 0);
  assign w750[49] = |(datain[115:112] ^ 1);
  assign w750[50] = |(datain[111:108] ^ 7);
  assign w750[51] = |(datain[107:104] ^ 3);
  assign w750[52] = |(datain[103:100] ^ 0);
  assign w750[53] = |(datain[99:96] ^ 3);
  assign w750[54] = |(datain[95:92] ^ 14);
  assign w750[55] = |(datain[91:88] ^ 9);
  assign w750[56] = |(datain[87:84] ^ 14);
  assign w750[57] = |(datain[83:80] ^ 5);
  assign w750[58] = |(datain[79:76] ^ 0);
  assign w750[59] = |(datain[75:72] ^ 0);
  assign w750[60] = |(datain[71:68] ^ 0);
  assign w750[61] = |(datain[67:64] ^ 5);
  assign w750[62] = |(datain[63:60] ^ 0);
  assign w750[63] = |(datain[59:56] ^ 2);
  assign w750[64] = |(datain[55:52] ^ 0);
  assign w750[65] = |(datain[51:48] ^ 0);
  assign w750[66] = |(datain[47:44] ^ 14);
  assign w750[67] = |(datain[43:40] ^ 8);
  assign w750[68] = |(datain[39:36] ^ 5);
  assign w750[69] = |(datain[35:32] ^ 13);
  assign w750[70] = |(datain[31:28] ^ 0);
  assign w750[71] = |(datain[27:24] ^ 1);
  assign w750[72] = |(datain[23:20] ^ 8);
  assign w750[73] = |(datain[19:16] ^ 11);
  assign comp[750] = ~(|w750);
  wire [38-1:0] w751;
  assign w751[0] = |(datain[311:308] ^ 0);
  assign w751[1] = |(datain[307:304] ^ 1);
  assign w751[2] = |(datain[303:300] ^ 11);
  assign w751[3] = |(datain[299:296] ^ 4);
  assign w751[4] = |(datain[295:292] ^ 4);
  assign w751[5] = |(datain[291:288] ^ 0);
  assign w751[6] = |(datain[287:284] ^ 12);
  assign w751[7] = |(datain[283:280] ^ 13);
  assign w751[8] = |(datain[279:276] ^ 2);
  assign w751[9] = |(datain[275:272] ^ 1);
  assign w751[10] = |(datain[271:268] ^ 7);
  assign w751[11] = |(datain[267:264] ^ 3);
  assign w751[12] = |(datain[263:260] ^ 0);
  assign w751[13] = |(datain[259:256] ^ 3);
  assign w751[14] = |(datain[255:252] ^ 14);
  assign w751[15] = |(datain[251:248] ^ 9);
  assign w751[16] = |(datain[247:244] ^ 4);
  assign w751[17] = |(datain[243:240] ^ 8);
  assign w751[18] = |(datain[239:236] ^ 0);
  assign w751[19] = |(datain[235:232] ^ 1);
  assign w751[20] = |(datain[231:228] ^ 2);
  assign w751[21] = |(datain[227:224] ^ 14);
  assign w751[22] = |(datain[223:220] ^ 8);
  assign w751[23] = |(datain[219:216] ^ 3);
  assign w751[24] = |(datain[215:212] ^ 2);
  assign w751[25] = |(datain[211:208] ^ 14);
  assign w751[26] = |(datain[207:204] ^ 1);
  assign w751[27] = |(datain[203:200] ^ 11);
  assign w751[28] = |(datain[199:196] ^ 0);
  assign w751[29] = |(datain[195:192] ^ 1);
  assign w751[30] = |(datain[191:188] ^ 0);
  assign w751[31] = |(datain[187:184] ^ 3);
  assign w751[32] = |(datain[183:180] ^ 3);
  assign w751[33] = |(datain[179:176] ^ 3);
  assign w751[34] = |(datain[175:172] ^ 12);
  assign w751[35] = |(datain[171:168] ^ 9);
  assign w751[36] = |(datain[167:164] ^ 3);
  assign w751[37] = |(datain[163:160] ^ 3);
  assign comp[751] = ~(|w751);
  wire [32-1:0] w752;
  assign w752[0] = |(datain[311:308] ^ 8);
  assign w752[1] = |(datain[307:304] ^ 3);
  assign w752[2] = |(datain[303:300] ^ 12);
  assign w752[3] = |(datain[299:296] ^ 7);
  assign w752[4] = |(datain[295:292] ^ 0);
  assign w752[5] = |(datain[291:288] ^ 7);
  assign w752[6] = |(datain[287:284] ^ 11);
  assign w752[7] = |(datain[283:280] ^ 9);
  assign w752[8] = |(datain[279:276] ^ 15);
  assign w752[9] = |(datain[275:272] ^ 9);
  assign w752[10] = |(datain[271:268] ^ 0);
  assign w752[11] = |(datain[267:264] ^ 4);
  assign w752[12] = |(datain[263:260] ^ 2);
  assign w752[13] = |(datain[259:256] ^ 14);
  assign w752[14] = |(datain[255:252] ^ 8);
  assign w752[15] = |(datain[251:248] ^ 0);
  assign w752[16] = |(datain[247:244] ^ 2);
  assign w752[17] = |(datain[243:240] ^ 13);
  assign w752[18] = |(datain[239:236] ^ 9);
  assign w752[19] = |(datain[235:232] ^ 3);
  assign w752[20] = |(datain[231:228] ^ 4);
  assign w752[21] = |(datain[227:224] ^ 7);
  assign w752[22] = |(datain[223:220] ^ 14);
  assign w752[23] = |(datain[219:216] ^ 2);
  assign w752[24] = |(datain[215:212] ^ 15);
  assign w752[25] = |(datain[211:208] ^ 9);
  assign w752[26] = |(datain[207:204] ^ 14);
  assign w752[27] = |(datain[203:200] ^ 9);
  assign w752[28] = |(datain[199:196] ^ 13);
  assign w752[29] = |(datain[195:192] ^ 10);
  assign w752[30] = |(datain[191:188] ^ 15);
  assign w752[31] = |(datain[187:184] ^ 14);
  assign comp[752] = ~(|w752);
  wire [42-1:0] w753;
  assign w753[0] = |(datain[311:308] ^ 12);
  assign w753[1] = |(datain[307:304] ^ 13);
  assign w753[2] = |(datain[303:300] ^ 2);
  assign w753[3] = |(datain[299:296] ^ 1);
  assign w753[4] = |(datain[295:292] ^ 3);
  assign w753[5] = |(datain[291:288] ^ 13);
  assign w753[6] = |(datain[287:284] ^ 14);
  assign w753[7] = |(datain[283:280] ^ 14);
  assign w753[8] = |(datain[279:276] ^ 15);
  assign w753[9] = |(datain[275:272] ^ 15);
  assign w753[10] = |(datain[271:268] ^ 7);
  assign w753[11] = |(datain[267:264] ^ 5);
  assign w753[12] = |(datain[263:260] ^ 0);
  assign w753[13] = |(datain[259:256] ^ 3);
  assign w753[14] = |(datain[255:252] ^ 14);
  assign w753[15] = |(datain[251:248] ^ 9);
  assign w753[16] = |(datain[247:244] ^ 13);
  assign w753[17] = |(datain[243:240] ^ 13);
  assign w753[18] = |(datain[239:236] ^ 0);
  assign w753[19] = |(datain[235:232] ^ 0);
  assign w753[20] = |(datain[231:228] ^ 0);
  assign w753[21] = |(datain[227:224] ^ 6);
  assign w753[22] = |(datain[223:220] ^ 11);
  assign w753[23] = |(datain[219:216] ^ 8);
  assign w753[24] = |(datain[215:212] ^ 2);
  assign w753[25] = |(datain[211:208] ^ 1);
  assign w753[26] = |(datain[207:204] ^ 3);
  assign w753[27] = |(datain[203:200] ^ 5);
  assign w753[28] = |(datain[199:196] ^ 12);
  assign w753[29] = |(datain[195:192] ^ 13);
  assign w753[30] = |(datain[191:188] ^ 2);
  assign w753[31] = |(datain[187:184] ^ 1);
  assign w753[32] = |(datain[183:180] ^ 2);
  assign w753[33] = |(datain[179:176] ^ 14);
  assign w753[34] = |(datain[175:172] ^ 8);
  assign w753[35] = |(datain[171:168] ^ 9);
  assign w753[36] = |(datain[167:164] ^ 1);
  assign w753[37] = |(datain[163:160] ^ 12);
  assign w753[38] = |(datain[159:156] ^ 2);
  assign w753[39] = |(datain[155:152] ^ 14);
  assign w753[40] = |(datain[151:148] ^ 8);
  assign w753[41] = |(datain[147:144] ^ 12);
  assign comp[753] = ~(|w753);
  wire [74-1:0] w754;
  assign w754[0] = |(datain[311:308] ^ 8);
  assign w754[1] = |(datain[307:304] ^ 13);
  assign w754[2] = |(datain[303:300] ^ 1);
  assign w754[3] = |(datain[299:296] ^ 6);
  assign w754[4] = |(datain[295:292] ^ 5);
  assign w754[5] = |(datain[291:288] ^ 10);
  assign w754[6] = |(datain[287:284] ^ 0);
  assign w754[7] = |(datain[283:280] ^ 1);
  assign w754[8] = |(datain[279:276] ^ 11);
  assign w754[9] = |(datain[275:272] ^ 4);
  assign w754[10] = |(datain[271:268] ^ 4);
  assign w754[11] = |(datain[267:264] ^ 0);
  assign w754[12] = |(datain[263:260] ^ 12);
  assign w754[13] = |(datain[259:256] ^ 13);
  assign w754[14] = |(datain[255:252] ^ 2);
  assign w754[15] = |(datain[251:248] ^ 1);
  assign w754[16] = |(datain[247:244] ^ 7);
  assign w754[17] = |(datain[243:240] ^ 2);
  assign w754[18] = |(datain[239:236] ^ 1);
  assign w754[19] = |(datain[235:232] ^ 0);
  assign w754[20] = |(datain[231:228] ^ 14);
  assign w754[21] = |(datain[227:224] ^ 8);
  assign w754[22] = |(datain[223:220] ^ 6);
  assign w754[23] = |(datain[219:216] ^ 8);
  assign w754[24] = |(datain[215:212] ^ 0);
  assign w754[25] = |(datain[211:208] ^ 1);
  assign w754[26] = |(datain[207:204] ^ 7);
  assign w754[27] = |(datain[203:200] ^ 2);
  assign w754[28] = |(datain[199:196] ^ 0);
  assign w754[29] = |(datain[195:192] ^ 11);
  assign w754[30] = |(datain[191:188] ^ 11);
  assign w754[31] = |(datain[187:184] ^ 9);
  assign w754[32] = |(datain[183:180] ^ 5);
  assign w754[33] = |(datain[179:176] ^ 2);
  assign w754[34] = |(datain[175:172] ^ 0);
  assign w754[35] = |(datain[171:168] ^ 7);
  assign w754[36] = |(datain[167:164] ^ 8);
  assign w754[37] = |(datain[163:160] ^ 13);
  assign w754[38] = |(datain[159:156] ^ 1);
  assign w754[39] = |(datain[155:152] ^ 6);
  assign w754[40] = |(datain[151:148] ^ 0);
  assign w754[41] = |(datain[147:144] ^ 0);
  assign w754[42] = |(datain[143:140] ^ 0);
  assign w754[43] = |(datain[139:136] ^ 1);
  assign w754[44] = |(datain[135:132] ^ 11);
  assign w754[45] = |(datain[131:128] ^ 4);
  assign w754[46] = |(datain[127:124] ^ 4);
  assign w754[47] = |(datain[123:120] ^ 0);
  assign w754[48] = |(datain[119:116] ^ 12);
  assign w754[49] = |(datain[115:112] ^ 13);
  assign w754[50] = |(datain[111:108] ^ 2);
  assign w754[51] = |(datain[107:104] ^ 1);
  assign w754[52] = |(datain[103:100] ^ 2);
  assign w754[53] = |(datain[99:96] ^ 14);
  assign w754[54] = |(datain[95:92] ^ 8);
  assign w754[55] = |(datain[91:88] ^ 11);
  assign w754[56] = |(datain[87:84] ^ 1);
  assign w754[57] = |(datain[83:80] ^ 14);
  assign w754[58] = |(datain[79:76] ^ 5);
  assign w754[59] = |(datain[75:72] ^ 2);
  assign w754[60] = |(datain[71:68] ^ 0);
  assign w754[61] = |(datain[67:64] ^ 1);
  assign w754[62] = |(datain[63:60] ^ 2);
  assign w754[63] = |(datain[59:56] ^ 14);
  assign w754[64] = |(datain[55:52] ^ 8);
  assign w754[65] = |(datain[51:48] ^ 11);
  assign w754[66] = |(datain[47:44] ^ 1);
  assign w754[67] = |(datain[43:40] ^ 6);
  assign w754[68] = |(datain[39:36] ^ 4);
  assign w754[69] = |(datain[35:32] ^ 10);
  assign w754[70] = |(datain[31:28] ^ 0);
  assign w754[71] = |(datain[27:24] ^ 1);
  assign w754[72] = |(datain[23:20] ^ 2);
  assign w754[73] = |(datain[19:16] ^ 14);
  assign comp[754] = ~(|w754);
  wire [46-1:0] w755;
  assign w755[0] = |(datain[311:308] ^ 1);
  assign w755[1] = |(datain[307:304] ^ 0);
  assign w755[2] = |(datain[303:300] ^ 0);
  assign w755[3] = |(datain[299:296] ^ 0);
  assign w755[4] = |(datain[295:292] ^ 2);
  assign w755[5] = |(datain[291:288] ^ 14);
  assign w755[6] = |(datain[287:284] ^ 0);
  assign w755[7] = |(datain[283:280] ^ 1);
  assign w755[8] = |(datain[279:276] ^ 4);
  assign w755[9] = |(datain[275:272] ^ 4);
  assign w755[10] = |(datain[271:268] ^ 7);
  assign w755[11] = |(datain[267:264] ^ 3);
  assign w755[12] = |(datain[263:260] ^ 2);
  assign w755[13] = |(datain[259:256] ^ 14);
  assign w755[14] = |(datain[255:252] ^ 8);
  assign w755[15] = |(datain[251:248] ^ 14);
  assign w755[16] = |(datain[247:244] ^ 5);
  assign w755[17] = |(datain[243:240] ^ 4);
  assign w755[18] = |(datain[239:236] ^ 7);
  assign w755[19] = |(datain[235:232] ^ 3);
  assign w755[20] = |(datain[231:228] ^ 3);
  assign w755[21] = |(datain[227:224] ^ 3);
  assign w755[22] = |(datain[223:220] ^ 12);
  assign w755[23] = |(datain[219:216] ^ 0);
  assign w755[24] = |(datain[215:212] ^ 2);
  assign w755[25] = |(datain[211:208] ^ 14);
  assign w755[26] = |(datain[207:204] ^ 8);
  assign w755[27] = |(datain[203:200] ^ 3);
  assign w755[28] = |(datain[199:196] ^ 4);
  assign w755[29] = |(datain[195:192] ^ 4);
  assign w755[30] = |(datain[191:188] ^ 3);
  assign w755[31] = |(datain[187:184] ^ 9);
  assign w755[32] = |(datain[183:180] ^ 1);
  assign w755[33] = |(datain[179:176] ^ 0);
  assign w755[34] = |(datain[175:172] ^ 2);
  assign w755[35] = |(datain[171:168] ^ 14);
  assign w755[36] = |(datain[167:164] ^ 15);
  assign w755[37] = |(datain[163:160] ^ 15);
  assign w755[38] = |(datain[159:156] ^ 6);
  assign w755[39] = |(datain[155:152] ^ 12);
  assign w755[40] = |(datain[151:148] ^ 3);
  assign w755[41] = |(datain[147:144] ^ 7);
  assign w755[42] = |(datain[143:140] ^ 5);
  assign w755[43] = |(datain[139:136] ^ 3);
  assign w755[44] = |(datain[135:132] ^ 4);
  assign w755[45] = |(datain[131:128] ^ 15);
  assign comp[755] = ~(|w755);
  wire [44-1:0] w756;
  assign w756[0] = |(datain[311:308] ^ 4);
  assign w756[1] = |(datain[307:304] ^ 11);
  assign w756[2] = |(datain[303:300] ^ 7);
  assign w756[3] = |(datain[299:296] ^ 4);
  assign w756[4] = |(datain[295:292] ^ 0);
  assign w756[5] = |(datain[291:288] ^ 3);
  assign w756[6] = |(datain[287:284] ^ 14);
  assign w756[7] = |(datain[283:280] ^ 9);
  assign w756[8] = |(datain[279:276] ^ 13);
  assign w756[9] = |(datain[275:272] ^ 11);
  assign w756[10] = |(datain[271:268] ^ 0);
  assign w756[11] = |(datain[267:264] ^ 2);
  assign w756[12] = |(datain[263:260] ^ 5);
  assign w756[13] = |(datain[259:256] ^ 0);
  assign w756[14] = |(datain[255:252] ^ 5);
  assign w756[15] = |(datain[251:248] ^ 3);
  assign w756[16] = |(datain[247:244] ^ 5);
  assign w756[17] = |(datain[243:240] ^ 1);
  assign w756[18] = |(datain[239:236] ^ 5);
  assign w756[19] = |(datain[235:232] ^ 2);
  assign w756[20] = |(datain[231:228] ^ 1);
  assign w756[21] = |(datain[227:224] ^ 14);
  assign w756[22] = |(datain[223:220] ^ 0);
  assign w756[23] = |(datain[219:216] ^ 6);
  assign w756[24] = |(datain[215:212] ^ 5);
  assign w756[25] = |(datain[211:208] ^ 6);
  assign w756[26] = |(datain[207:204] ^ 5);
  assign w756[27] = |(datain[203:200] ^ 7);
  assign w756[28] = |(datain[199:196] ^ 2);
  assign w756[29] = |(datain[195:192] ^ 14);
  assign w756[30] = |(datain[191:188] ^ 8);
  assign w756[31] = |(datain[187:184] ^ 9);
  assign w756[32] = |(datain[183:180] ^ 1);
  assign w756[33] = |(datain[179:176] ^ 6);
  assign w756[34] = |(datain[175:172] ^ 4);
  assign w756[35] = |(datain[171:168] ^ 14);
  assign w756[36] = |(datain[167:164] ^ 0);
  assign w756[37] = |(datain[163:160] ^ 1);
  assign w756[38] = |(datain[159:156] ^ 2);
  assign w756[39] = |(datain[155:152] ^ 14);
  assign w756[40] = |(datain[151:148] ^ 8);
  assign w756[41] = |(datain[147:144] ^ 12);
  assign w756[42] = |(datain[143:140] ^ 1);
  assign w756[43] = |(datain[139:136] ^ 14);
  assign comp[756] = ~(|w756);
  wire [42-1:0] w757;
  assign w757[0] = |(datain[311:308] ^ 7);
  assign w757[1] = |(datain[307:304] ^ 4);
  assign w757[2] = |(datain[303:300] ^ 0);
  assign w757[3] = |(datain[299:296] ^ 3);
  assign w757[4] = |(datain[295:292] ^ 14);
  assign w757[5] = |(datain[291:288] ^ 9);
  assign w757[6] = |(datain[287:284] ^ 11);
  assign w757[7] = |(datain[283:280] ^ 10);
  assign w757[8] = |(datain[279:276] ^ 0);
  assign w757[9] = |(datain[275:272] ^ 1);
  assign w757[10] = |(datain[271:268] ^ 5);
  assign w757[11] = |(datain[267:264] ^ 0);
  assign w757[12] = |(datain[263:260] ^ 5);
  assign w757[13] = |(datain[259:256] ^ 3);
  assign w757[14] = |(datain[255:252] ^ 5);
  assign w757[15] = |(datain[251:248] ^ 1);
  assign w757[16] = |(datain[247:244] ^ 5);
  assign w757[17] = |(datain[243:240] ^ 2);
  assign w757[18] = |(datain[239:236] ^ 1);
  assign w757[19] = |(datain[235:232] ^ 14);
  assign w757[20] = |(datain[231:228] ^ 0);
  assign w757[21] = |(datain[227:224] ^ 6);
  assign w757[22] = |(datain[223:220] ^ 5);
  assign w757[23] = |(datain[219:216] ^ 6);
  assign w757[24] = |(datain[215:212] ^ 5);
  assign w757[25] = |(datain[211:208] ^ 7);
  assign w757[26] = |(datain[207:204] ^ 2);
  assign w757[27] = |(datain[203:200] ^ 14);
  assign w757[28] = |(datain[199:196] ^ 8);
  assign w757[29] = |(datain[195:192] ^ 9);
  assign w757[30] = |(datain[191:188] ^ 1);
  assign w757[31] = |(datain[187:184] ^ 6);
  assign w757[32] = |(datain[183:180] ^ 4);
  assign w757[33] = |(datain[179:176] ^ 7);
  assign w757[34] = |(datain[175:172] ^ 0);
  assign w757[35] = |(datain[171:168] ^ 1);
  assign w757[36] = |(datain[167:164] ^ 2);
  assign w757[37] = |(datain[163:160] ^ 14);
  assign w757[38] = |(datain[159:156] ^ 8);
  assign w757[39] = |(datain[155:152] ^ 12);
  assign w757[40] = |(datain[151:148] ^ 1);
  assign w757[41] = |(datain[147:144] ^ 14);
  assign comp[757] = ~(|w757);
  wire [74-1:0] w758;
  assign w758[0] = |(datain[311:308] ^ 1);
  assign w758[1] = |(datain[307:304] ^ 15);
  assign w758[2] = |(datain[303:300] ^ 8);
  assign w758[3] = |(datain[299:296] ^ 11);
  assign w758[4] = |(datain[295:292] ^ 13);
  assign w758[5] = |(datain[291:288] ^ 3);
  assign w758[6] = |(datain[287:284] ^ 15);
  assign w758[7] = |(datain[283:280] ^ 2);
  assign w758[8] = |(datain[279:276] ^ 12);
  assign w758[9] = |(datain[275:272] ^ 1);
  assign w758[10] = |(datain[271:268] ^ 11);
  assign w758[11] = |(datain[267:264] ^ 4);
  assign w758[12] = |(datain[263:260] ^ 4);
  assign w758[13] = |(datain[259:256] ^ 0);
  assign w758[14] = |(datain[255:252] ^ 12);
  assign w758[15] = |(datain[251:248] ^ 13);
  assign w758[16] = |(datain[247:244] ^ 2);
  assign w758[17] = |(datain[243:240] ^ 1);
  assign w758[18] = |(datain[239:236] ^ 11);
  assign w758[19] = |(datain[235:232] ^ 8);
  assign w758[20] = |(datain[231:228] ^ 1);
  assign w758[21] = |(datain[227:224] ^ 7);
  assign w758[22] = |(datain[223:220] ^ 15);
  assign w758[23] = |(datain[219:216] ^ 15);
  assign w758[24] = |(datain[215:212] ^ 11);
  assign w758[25] = |(datain[211:208] ^ 10);
  assign w758[26] = |(datain[207:204] ^ 3);
  assign w758[27] = |(datain[203:200] ^ 8);
  assign w758[28] = |(datain[199:196] ^ 0);
  assign w758[29] = |(datain[195:192] ^ 0);
  assign w758[30] = |(datain[191:188] ^ 11);
  assign w758[31] = |(datain[187:184] ^ 9);
  assign w758[32] = |(datain[183:180] ^ 3);
  assign w758[33] = |(datain[179:176] ^ 6);
  assign w758[34] = |(datain[175:172] ^ 4);
  assign w758[35] = |(datain[171:168] ^ 1);
  assign w758[36] = |(datain[167:164] ^ 15);
  assign w758[37] = |(datain[163:160] ^ 4);
  assign w758[38] = |(datain[159:156] ^ 1);
  assign w758[39] = |(datain[155:152] ^ 15);
  assign w758[40] = |(datain[151:148] ^ 12);
  assign w758[41] = |(datain[147:144] ^ 6);
  assign w758[42] = |(datain[143:140] ^ 0);
  assign w758[43] = |(datain[139:136] ^ 6);
  assign w758[44] = |(datain[135:132] ^ 0);
  assign w758[45] = |(datain[131:128] ^ 4);
  assign w758[46] = |(datain[127:124] ^ 0);
  assign w758[47] = |(datain[123:120] ^ 0);
  assign w758[48] = |(datain[119:116] ^ 0);
  assign w758[49] = |(datain[115:112] ^ 0);
  assign w758[50] = |(datain[111:108] ^ 15);
  assign w758[51] = |(datain[107:104] ^ 15);
  assign w758[52] = |(datain[103:100] ^ 1);
  assign w758[53] = |(datain[99:96] ^ 11);
  assign w758[54] = |(datain[95:92] ^ 14);
  assign w758[55] = |(datain[91:88] ^ 11);
  assign w758[56] = |(datain[87:84] ^ 1);
  assign w758[57] = |(datain[83:80] ^ 12);
  assign w758[58] = |(datain[79:76] ^ 9);
  assign w758[59] = |(datain[75:72] ^ 0);
  assign w758[60] = |(datain[71:68] ^ 1);
  assign w758[61] = |(datain[67:64] ^ 15);
  assign w758[62] = |(datain[63:60] ^ 12);
  assign w758[63] = |(datain[59:56] ^ 13);
  assign w758[64] = |(datain[55:52] ^ 1);
  assign w758[65] = |(datain[51:48] ^ 1);
  assign w758[66] = |(datain[47:44] ^ 2);
  assign w758[67] = |(datain[43:40] ^ 4);
  assign w758[68] = |(datain[39:36] ^ 0);
  assign w758[69] = |(datain[35:32] ^ 2);
  assign w758[70] = |(datain[31:28] ^ 13);
  assign w758[71] = |(datain[27:24] ^ 0);
  assign w758[72] = |(datain[23:20] ^ 14);
  assign w758[73] = |(datain[19:16] ^ 8);
  assign comp[758] = ~(|w758);
  wire [32-1:0] w759;
  assign w759[0] = |(datain[311:308] ^ 12);
  assign w759[1] = |(datain[307:304] ^ 13);
  assign w759[2] = |(datain[303:300] ^ 2);
  assign w759[3] = |(datain[299:296] ^ 1);
  assign w759[4] = |(datain[295:292] ^ 8);
  assign w759[5] = |(datain[291:288] ^ 11);
  assign w759[6] = |(datain[287:284] ^ 13);
  assign w759[7] = |(datain[283:280] ^ 5);
  assign w759[8] = |(datain[279:276] ^ 8);
  assign w759[9] = |(datain[275:272] ^ 1);
  assign w759[10] = |(datain[271:268] ^ 12);
  assign w759[11] = |(datain[267:264] ^ 2);
  assign w759[12] = |(datain[263:260] ^ 5);
  assign w759[13] = |(datain[259:256] ^ 4);
  assign w759[14] = |(datain[255:252] ^ 0);
  assign w759[15] = |(datain[251:248] ^ 2);
  assign w759[16] = |(datain[247:244] ^ 11);
  assign w759[17] = |(datain[243:240] ^ 9);
  assign w759[18] = |(datain[239:236] ^ 0);
  assign w759[19] = |(datain[235:232] ^ 7);
  assign w759[20] = |(datain[231:228] ^ 0);
  assign w759[21] = |(datain[227:224] ^ 0);
  assign w759[22] = |(datain[223:220] ^ 11);
  assign w759[23] = |(datain[219:216] ^ 4);
  assign w759[24] = |(datain[215:212] ^ 3);
  assign w759[25] = |(datain[211:208] ^ 15);
  assign w759[26] = |(datain[207:204] ^ 12);
  assign w759[27] = |(datain[203:200] ^ 13);
  assign w759[28] = |(datain[199:196] ^ 2);
  assign w759[29] = |(datain[195:192] ^ 1);
  assign w759[30] = |(datain[191:188] ^ 15);
  assign w759[31] = |(datain[187:184] ^ 12);
  assign comp[759] = ~(|w759);
  wire [42-1:0] w760;
  assign w760[0] = |(datain[311:308] ^ 11);
  assign w760[1] = |(datain[307:304] ^ 14);
  assign w760[2] = |(datain[303:300] ^ 1);
  assign w760[3] = |(datain[299:296] ^ 3);
  assign w760[4] = |(datain[295:292] ^ 0);
  assign w760[5] = |(datain[291:288] ^ 5);
  assign w760[6] = |(datain[287:284] ^ 8);
  assign w760[7] = |(datain[283:280] ^ 11);
  assign w760[8] = |(datain[279:276] ^ 15);
  assign w760[9] = |(datain[275:272] ^ 14);
  assign w760[10] = |(datain[271:268] ^ 8);
  assign w760[11] = |(datain[267:264] ^ 1);
  assign w760[12] = |(datain[263:260] ^ 12);
  assign w760[13] = |(datain[259:256] ^ 7);
  assign w760[14] = |(datain[255:252] ^ 6);
  assign w760[15] = |(datain[251:248] ^ 3);
  assign w760[16] = |(datain[247:244] ^ 0);
  assign w760[17] = |(datain[243:240] ^ 2);
  assign w760[18] = |(datain[239:236] ^ 9);
  assign w760[19] = |(datain[235:232] ^ 11);
  assign w760[20] = |(datain[231:228] ^ 13);
  assign w760[21] = |(datain[227:224] ^ 11);
  assign w760[22] = |(datain[223:220] ^ 14);
  assign w760[23] = |(datain[219:216] ^ 3);
  assign w760[24] = |(datain[215:212] ^ 9);
  assign w760[25] = |(datain[211:208] ^ 11);
  assign w760[26] = |(datain[207:204] ^ 2);
  assign w760[27] = |(datain[203:200] ^ 14);
  assign w760[28] = |(datain[199:196] ^ 13);
  assign w760[29] = |(datain[195:192] ^ 13);
  assign w760[30] = |(datain[191:188] ^ 0);
  assign w760[31] = |(datain[187:184] ^ 5);
  assign w760[32] = |(datain[183:180] ^ 9);
  assign w760[33] = |(datain[179:176] ^ 11);
  assign w760[34] = |(datain[175:172] ^ 2);
  assign w760[35] = |(datain[171:168] ^ 14);
  assign w760[36] = |(datain[167:164] ^ 13);
  assign w760[37] = |(datain[163:160] ^ 13);
  assign w760[38] = |(datain[159:156] ^ 1);
  assign w760[39] = |(datain[155:152] ^ 5);
  assign w760[40] = |(datain[151:148] ^ 9);
  assign w760[41] = |(datain[147:144] ^ 11);
  assign comp[760] = ~(|w760);
  wire [44-1:0] w761;
  assign w761[0] = |(datain[311:308] ^ 10);
  assign w761[1] = |(datain[307:304] ^ 3);
  assign w761[2] = |(datain[303:300] ^ 6);
  assign w761[3] = |(datain[299:296] ^ 0);
  assign w761[4] = |(datain[295:292] ^ 0);
  assign w761[5] = |(datain[291:288] ^ 0);
  assign w761[6] = |(datain[287:284] ^ 8);
  assign w761[7] = |(datain[283:280] ^ 12);
  assign w761[8] = |(datain[279:276] ^ 0);
  assign w761[9] = |(datain[275:272] ^ 6);
  assign w761[10] = |(datain[271:268] ^ 6);
  assign w761[11] = |(datain[267:264] ^ 2);
  assign w761[12] = |(datain[263:260] ^ 0);
  assign w761[13] = |(datain[259:256] ^ 0);
  assign w761[14] = |(datain[255:252] ^ 12);
  assign w761[15] = |(datain[251:248] ^ 7);
  assign w761[16] = |(datain[247:244] ^ 0);
  assign w761[17] = |(datain[243:240] ^ 6);
  assign w761[18] = |(datain[239:236] ^ 4);
  assign w761[19] = |(datain[235:232] ^ 12);
  assign w761[20] = |(datain[231:228] ^ 0);
  assign w761[21] = |(datain[227:224] ^ 0);
  assign w761[22] = |(datain[223:220] ^ 7);
  assign w761[23] = |(datain[219:216] ^ 15);
  assign w761[24] = |(datain[215:212] ^ 7);
  assign w761[25] = |(datain[211:208] ^ 12);
  assign w761[26] = |(datain[207:204] ^ 8);
  assign w761[27] = |(datain[203:200] ^ 12);
  assign w761[28] = |(datain[199:196] ^ 0);
  assign w761[29] = |(datain[195:192] ^ 14);
  assign w761[30] = |(datain[191:188] ^ 4);
  assign w761[31] = |(datain[187:184] ^ 14);
  assign w761[32] = |(datain[183:180] ^ 0);
  assign w761[33] = |(datain[179:176] ^ 0);
  assign w761[34] = |(datain[175:172] ^ 12);
  assign w761[35] = |(datain[171:168] ^ 7);
  assign w761[36] = |(datain[167:164] ^ 0);
  assign w761[37] = |(datain[163:160] ^ 6);
  assign w761[38] = |(datain[159:156] ^ 7);
  assign w761[39] = |(datain[155:152] ^ 0);
  assign w761[40] = |(datain[151:148] ^ 0);
  assign w761[41] = |(datain[147:144] ^ 0);
  assign w761[42] = |(datain[143:140] ^ 4);
  assign w761[43] = |(datain[139:136] ^ 13);
  assign comp[761] = ~(|w761);
  wire [42-1:0] w762;
  assign w762[0] = |(datain[311:308] ^ 5);
  assign w762[1] = |(datain[307:304] ^ 14);
  assign w762[2] = |(datain[303:300] ^ 8);
  assign w762[3] = |(datain[299:296] ^ 1);
  assign w762[4] = |(datain[295:292] ^ 14);
  assign w762[5] = |(datain[291:288] ^ 14);
  assign w762[6] = |(datain[287:284] ^ 4);
  assign w762[7] = |(datain[283:280] ^ 3);
  assign w762[8] = |(datain[279:276] ^ 0);
  assign w762[9] = |(datain[275:272] ^ 6);
  assign w762[10] = |(datain[271:268] ^ 8);
  assign w762[11] = |(datain[267:264] ^ 11);
  assign w762[12] = |(datain[263:260] ^ 15);
  assign w762[13] = |(datain[259:256] ^ 14);
  assign w762[14] = |(datain[255:252] ^ 5);
  assign w762[15] = |(datain[251:248] ^ 7);
  assign w762[16] = |(datain[247:244] ^ 5);
  assign w762[17] = |(datain[243:240] ^ 0);
  assign w762[18] = |(datain[239:236] ^ 1);
  assign w762[19] = |(datain[235:232] ^ 14);
  assign w762[20] = |(datain[231:228] ^ 0);
  assign w762[21] = |(datain[227:224] ^ 6);
  assign w762[22] = |(datain[223:220] ^ 0);
  assign w762[23] = |(datain[219:216] ^ 14);
  assign w762[24] = |(datain[215:212] ^ 0);
  assign w762[25] = |(datain[211:208] ^ 7);
  assign w762[26] = |(datain[207:204] ^ 0);
  assign w762[27] = |(datain[203:200] ^ 14);
  assign w762[28] = |(datain[199:196] ^ 1);
  assign w762[29] = |(datain[195:192] ^ 15);
  assign w762[30] = |(datain[191:188] ^ 11);
  assign w762[31] = |(datain[187:184] ^ 6);
  assign w762[32] = |(datain[183:180] ^ 5);
  assign w762[33] = |(datain[179:176] ^ 8);
  assign w762[34] = |(datain[175:172] ^ 11);
  assign w762[35] = |(datain[171:168] ^ 9);
  assign w762[36] = |(datain[167:164] ^ 4);
  assign w762[37] = |(datain[163:160] ^ 0);
  assign w762[38] = |(datain[159:156] ^ 0);
  assign w762[39] = |(datain[155:152] ^ 6);
  assign w762[40] = |(datain[151:148] ^ 10);
  assign w762[41] = |(datain[147:144] ^ 12);
  assign comp[762] = ~(|w762);
  wire [74-1:0] w763;
  assign w763[0] = |(datain[311:308] ^ 2);
  assign w763[1] = |(datain[307:304] ^ 7);
  assign w763[2] = |(datain[303:300] ^ 12);
  assign w763[3] = |(datain[299:296] ^ 14);
  assign w763[4] = |(datain[295:292] ^ 1);
  assign w763[5] = |(datain[291:288] ^ 13);
  assign w763[6] = |(datain[287:284] ^ 3);
  assign w763[7] = |(datain[283:280] ^ 12);
  assign w763[8] = |(datain[279:276] ^ 11);
  assign w763[9] = |(datain[275:272] ^ 9);
  assign w763[10] = |(datain[271:268] ^ 9);
  assign w763[11] = |(datain[267:264] ^ 9);
  assign w763[12] = |(datain[263:260] ^ 9);
  assign w763[13] = |(datain[259:256] ^ 10);
  assign w763[14] = |(datain[255:252] ^ 5);
  assign w763[15] = |(datain[251:248] ^ 7);
  assign w763[16] = |(datain[247:244] ^ 7);
  assign w763[17] = |(datain[243:240] ^ 3);
  assign w763[18] = |(datain[239:236] ^ 9);
  assign w763[19] = |(datain[235:232] ^ 5);
  assign w763[20] = |(datain[231:228] ^ 1);
  assign w763[21] = |(datain[227:224] ^ 10);
  assign w763[22] = |(datain[223:220] ^ 5);
  assign w763[23] = |(datain[219:216] ^ 6);
  assign w763[24] = |(datain[215:212] ^ 7);
  assign w763[25] = |(datain[211:208] ^ 10);
  assign w763[26] = |(datain[207:204] ^ 3);
  assign w763[27] = |(datain[203:200] ^ 8);
  assign w763[28] = |(datain[199:196] ^ 2);
  assign w763[29] = |(datain[195:192] ^ 11);
  assign w763[30] = |(datain[191:188] ^ 2);
  assign w763[31] = |(datain[187:184] ^ 6);
  assign w763[32] = |(datain[183:180] ^ 3);
  assign w763[33] = |(datain[179:176] ^ 13);
  assign w763[34] = |(datain[175:172] ^ 2);
  assign w763[35] = |(datain[171:168] ^ 4);
  assign w763[36] = |(datain[167:164] ^ 4);
  assign w763[37] = |(datain[163:160] ^ 8);
  assign w763[38] = |(datain[159:156] ^ 6);
  assign w763[39] = |(datain[155:152] ^ 2);
  assign w763[40] = |(datain[151:148] ^ 6);
  assign w763[41] = |(datain[147:144] ^ 6);
  assign w763[42] = |(datain[143:140] ^ 2);
  assign w763[43] = |(datain[139:136] ^ 11);
  assign w763[44] = |(datain[135:132] ^ 2);
  assign w763[45] = |(datain[131:128] ^ 7);
  assign w763[46] = |(datain[127:124] ^ 2);
  assign w763[47] = |(datain[123:120] ^ 5);
  assign w763[48] = |(datain[119:116] ^ 14);
  assign w763[49] = |(datain[115:112] ^ 0);
  assign w763[50] = |(datain[111:108] ^ 6);
  assign w763[51] = |(datain[107:104] ^ 0);
  assign w763[52] = |(datain[103:100] ^ 3);
  assign w763[53] = |(datain[99:96] ^ 4);
  assign w763[54] = |(datain[95:92] ^ 0);
  assign w763[55] = |(datain[91:88] ^ 11);
  assign w763[56] = |(datain[87:84] ^ 6);
  assign w763[57] = |(datain[83:80] ^ 7);
  assign w763[58] = |(datain[79:76] ^ 0);
  assign w763[59] = |(datain[75:72] ^ 4);
  assign w763[60] = |(datain[71:68] ^ 4);
  assign w763[61] = |(datain[67:64] ^ 2);
  assign w763[62] = |(datain[63:60] ^ 9);
  assign w763[63] = |(datain[59:56] ^ 1);
  assign w763[64] = |(datain[55:52] ^ 7);
  assign w763[65] = |(datain[51:48] ^ 14);
  assign w763[66] = |(datain[47:44] ^ 2);
  assign w763[67] = |(datain[43:40] ^ 12);
  assign w763[68] = |(datain[39:36] ^ 3);
  assign w763[69] = |(datain[35:32] ^ 9);
  assign w763[70] = |(datain[31:28] ^ 7);
  assign w763[71] = |(datain[27:24] ^ 0);
  assign w763[72] = |(datain[23:20] ^ 9);
  assign w763[73] = |(datain[19:16] ^ 9);
  assign comp[763] = ~(|w763);
  wire [74-1:0] w764;
  assign w764[0] = |(datain[311:308] ^ 0);
  assign w764[1] = |(datain[307:304] ^ 13);
  assign w764[2] = |(datain[303:300] ^ 0);
  assign w764[3] = |(datain[299:296] ^ 10);
  assign w764[4] = |(datain[295:292] ^ 6);
  assign w764[5] = |(datain[291:288] ^ 6);
  assign w764[6] = |(datain[287:284] ^ 6);
  assign w764[7] = |(datain[283:280] ^ 15);
  assign w764[8] = |(datain[279:276] ^ 7);
  assign w764[9] = |(datain[275:272] ^ 2);
  assign w764[10] = |(datain[271:268] ^ 2);
  assign w764[11] = |(datain[267:264] ^ 0);
  assign w764[12] = |(datain[263:260] ^ 2);
  assign w764[13] = |(datain[259:256] ^ 5);
  assign w764[14] = |(datain[255:252] ^ 2);
  assign w764[15] = |(datain[251:248] ^ 5);
  assign w764[16] = |(datain[247:244] ^ 6);
  assign w764[17] = |(datain[243:240] ^ 2);
  assign w764[18] = |(datain[239:236] ^ 2);
  assign w764[19] = |(datain[235:232] ^ 0);
  assign w764[20] = |(datain[231:228] ^ 6);
  assign w764[21] = |(datain[227:224] ^ 9);
  assign w764[22] = |(datain[223:220] ^ 6);
  assign w764[23] = |(datain[219:216] ^ 14);
  assign w764[24] = |(datain[215:212] ^ 2);
  assign w764[25] = |(datain[211:208] ^ 0);
  assign w764[26] = |(datain[207:204] ^ 2);
  assign w764[27] = |(datain[203:200] ^ 8);
  assign w764[28] = |(datain[199:196] ^ 2);
  assign w764[29] = |(datain[195:192] ^ 10);
  assign w764[30] = |(datain[191:188] ^ 2);
  assign w764[31] = |(datain[187:184] ^ 14);
  assign w764[32] = |(datain[183:180] ^ 6);
  assign w764[33] = |(datain[179:176] ^ 2);
  assign w764[34] = |(datain[175:172] ^ 6);
  assign w764[35] = |(datain[171:168] ^ 1);
  assign w764[36] = |(datain[167:164] ^ 7);
  assign w764[37] = |(datain[163:160] ^ 4);
  assign w764[38] = |(datain[159:156] ^ 2);
  assign w764[39] = |(datain[155:152] ^ 9);
  assign w764[40] = |(datain[151:148] ^ 2);
  assign w764[41] = |(datain[147:144] ^ 0);
  assign w764[42] = |(datain[143:140] ^ 6);
  assign w764[43] = |(datain[139:136] ^ 4);
  assign w764[44] = |(datain[135:132] ^ 6);
  assign w764[45] = |(datain[131:128] ^ 15);
  assign w764[46] = |(datain[127:124] ^ 2);
  assign w764[47] = |(datain[123:120] ^ 0);
  assign w764[48] = |(datain[119:116] ^ 6);
  assign w764[49] = |(datain[115:112] ^ 3);
  assign w764[50] = |(datain[111:108] ^ 6);
  assign w764[51] = |(datain[107:104] ^ 1);
  assign w764[52] = |(datain[103:100] ^ 6);
  assign w764[53] = |(datain[99:96] ^ 12);
  assign w764[54] = |(datain[95:92] ^ 6);
  assign w764[55] = |(datain[91:88] ^ 12);
  assign w764[56] = |(datain[87:84] ^ 2);
  assign w764[57] = |(datain[83:80] ^ 0);
  assign w764[58] = |(datain[79:76] ^ 2);
  assign w764[59] = |(datain[75:72] ^ 5);
  assign w764[60] = |(datain[71:68] ^ 3);
  assign w764[61] = |(datain[67:64] ^ 0);
  assign w764[62] = |(datain[63:60] ^ 2);
  assign w764[63] = |(datain[59:56] ^ 0);
  assign w764[64] = |(datain[55:52] ^ 3);
  assign w764[65] = |(datain[51:48] ^ 4);
  assign w764[66] = |(datain[47:44] ^ 2);
  assign w764[67] = |(datain[43:40] ^ 0);
  assign w764[68] = |(datain[39:36] ^ 2);
  assign w764[69] = |(datain[35:32] ^ 5);
  assign w764[70] = |(datain[31:28] ^ 2);
  assign w764[71] = |(datain[27:24] ^ 5);
  assign w764[72] = |(datain[23:20] ^ 6);
  assign w764[73] = |(datain[19:16] ^ 2);
  assign comp[764] = ~(|w764);
  wire [74-1:0] w765;
  assign w765[0] = |(datain[311:308] ^ 0);
  assign w765[1] = |(datain[307:304] ^ 13);
  assign w765[2] = |(datain[303:300] ^ 0);
  assign w765[3] = |(datain[299:296] ^ 10);
  assign w765[4] = |(datain[295:292] ^ 6);
  assign w765[5] = |(datain[291:288] ^ 6);
  assign w765[6] = |(datain[287:284] ^ 6);
  assign w765[7] = |(datain[283:280] ^ 15);
  assign w765[8] = |(datain[279:276] ^ 7);
  assign w765[9] = |(datain[275:272] ^ 2);
  assign w765[10] = |(datain[271:268] ^ 2);
  assign w765[11] = |(datain[267:264] ^ 0);
  assign w765[12] = |(datain[263:260] ^ 2);
  assign w765[13] = |(datain[259:256] ^ 5);
  assign w765[14] = |(datain[255:252] ^ 2);
  assign w765[15] = |(datain[251:248] ^ 5);
  assign w765[16] = |(datain[247:244] ^ 6);
  assign w765[17] = |(datain[243:240] ^ 6);
  assign w765[18] = |(datain[239:236] ^ 2);
  assign w765[19] = |(datain[235:232] ^ 0);
  assign w765[20] = |(datain[231:228] ^ 6);
  assign w765[21] = |(datain[227:224] ^ 9);
  assign w765[22] = |(datain[223:220] ^ 6);
  assign w765[23] = |(datain[219:216] ^ 14);
  assign w765[24] = |(datain[215:212] ^ 2);
  assign w765[25] = |(datain[211:208] ^ 0);
  assign w765[26] = |(datain[207:204] ^ 2);
  assign w765[27] = |(datain[203:200] ^ 8);
  assign w765[28] = |(datain[199:196] ^ 2);
  assign w765[29] = |(datain[195:192] ^ 10);
  assign w765[30] = |(datain[191:188] ^ 2);
  assign w765[31] = |(datain[187:184] ^ 14);
  assign w765[32] = |(datain[183:180] ^ 6);
  assign w765[33] = |(datain[179:176] ^ 2);
  assign w765[34] = |(datain[175:172] ^ 6);
  assign w765[35] = |(datain[171:168] ^ 1);
  assign w765[36] = |(datain[167:164] ^ 7);
  assign w765[37] = |(datain[163:160] ^ 4);
  assign w765[38] = |(datain[159:156] ^ 2);
  assign w765[39] = |(datain[155:152] ^ 9);
  assign w765[40] = |(datain[151:148] ^ 2);
  assign w765[41] = |(datain[147:144] ^ 0);
  assign w765[42] = |(datain[143:140] ^ 6);
  assign w765[43] = |(datain[139:136] ^ 4);
  assign w765[44] = |(datain[135:132] ^ 6);
  assign w765[45] = |(datain[131:128] ^ 15);
  assign w765[46] = |(datain[127:124] ^ 2);
  assign w765[47] = |(datain[123:120] ^ 0);
  assign w765[48] = |(datain[119:116] ^ 6);
  assign w765[49] = |(datain[115:112] ^ 3);
  assign w765[50] = |(datain[111:108] ^ 6);
  assign w765[51] = |(datain[107:104] ^ 1);
  assign w765[52] = |(datain[103:100] ^ 6);
  assign w765[53] = |(datain[99:96] ^ 12);
  assign w765[54] = |(datain[95:92] ^ 6);
  assign w765[55] = |(datain[91:88] ^ 12);
  assign w765[56] = |(datain[87:84] ^ 2);
  assign w765[57] = |(datain[83:80] ^ 0);
  assign w765[58] = |(datain[79:76] ^ 2);
  assign w765[59] = |(datain[75:72] ^ 5);
  assign w765[60] = |(datain[71:68] ^ 3);
  assign w765[61] = |(datain[67:64] ^ 0);
  assign w765[62] = |(datain[63:60] ^ 2);
  assign w765[63] = |(datain[59:56] ^ 0);
  assign w765[64] = |(datain[55:52] ^ 3);
  assign w765[65] = |(datain[51:48] ^ 7);
  assign w765[66] = |(datain[47:44] ^ 2);
  assign w765[67] = |(datain[43:40] ^ 0);
  assign w765[68] = |(datain[39:36] ^ 2);
  assign w765[69] = |(datain[35:32] ^ 5);
  assign w765[70] = |(datain[31:28] ^ 2);
  assign w765[71] = |(datain[27:24] ^ 5);
  assign w765[72] = |(datain[23:20] ^ 6);
  assign w765[73] = |(datain[19:16] ^ 6);
  assign comp[765] = ~(|w765);
  wire [76-1:0] w766;
  assign w766[0] = |(datain[311:308] ^ 3);
  assign w766[1] = |(datain[307:304] ^ 3);
  assign w766[2] = |(datain[303:300] ^ 12);
  assign w766[3] = |(datain[299:296] ^ 0);
  assign w766[4] = |(datain[295:292] ^ 9);
  assign w766[5] = |(datain[291:288] ^ 14);
  assign w766[6] = |(datain[287:284] ^ 9);
  assign w766[7] = |(datain[283:280] ^ 15);
  assign w766[8] = |(datain[279:276] ^ 8);
  assign w766[9] = |(datain[275:272] ^ 0);
  assign w766[10] = |(datain[271:268] ^ 12);
  assign w766[11] = |(datain[267:264] ^ 4);
  assign w766[12] = |(datain[263:260] ^ 3);
  assign w766[13] = |(datain[259:256] ^ 14);
  assign w766[14] = |(datain[255:252] ^ 5);
  assign w766[15] = |(datain[251:248] ^ 0);
  assign w766[16] = |(datain[247:244] ^ 8);
  assign w766[17] = |(datain[243:240] ^ 11);
  assign w766[18] = |(datain[239:236] ^ 0);
  assign w766[19] = |(datain[235:232] ^ 14);
  assign w766[20] = |(datain[231:228] ^ 3);
  assign w766[21] = |(datain[227:224] ^ 6);
  assign w766[22] = |(datain[223:220] ^ 0);
  assign w766[23] = |(datain[219:216] ^ 1);
  assign w766[24] = |(datain[215:212] ^ 11);
  assign w766[25] = |(datain[211:208] ^ 10);
  assign w766[26] = |(datain[207:204] ^ 0);
  assign w766[27] = |(datain[203:200] ^ 0);
  assign w766[28] = |(datain[199:196] ^ 0);
  assign w766[29] = |(datain[195:192] ^ 1);
  assign w766[30] = |(datain[191:188] ^ 12);
  assign w766[31] = |(datain[187:184] ^ 13);
  assign w766[32] = |(datain[183:180] ^ 2);
  assign w766[33] = |(datain[179:176] ^ 1);
  assign w766[34] = |(datain[175:172] ^ 11);
  assign w766[35] = |(datain[171:168] ^ 8);
  assign w766[36] = |(datain[167:164] ^ 0);
  assign w766[37] = |(datain[163:160] ^ 2);
  assign w766[38] = |(datain[159:156] ^ 4);
  assign w766[39] = |(datain[155:152] ^ 2);
  assign w766[40] = |(datain[151:148] ^ 3);
  assign w766[41] = |(datain[147:144] ^ 3);
  assign w766[42] = |(datain[143:140] ^ 12);
  assign w766[43] = |(datain[139:136] ^ 9);
  assign w766[44] = |(datain[135:132] ^ 3);
  assign w766[45] = |(datain[131:128] ^ 3);
  assign w766[46] = |(datain[127:124] ^ 13);
  assign w766[47] = |(datain[123:120] ^ 2);
  assign w766[48] = |(datain[119:116] ^ 12);
  assign w766[49] = |(datain[115:112] ^ 13);
  assign w766[50] = |(datain[111:108] ^ 2);
  assign w766[51] = |(datain[107:104] ^ 1);
  assign w766[52] = |(datain[103:100] ^ 5);
  assign w766[53] = |(datain[99:96] ^ 8);
  assign w766[54] = |(datain[95:92] ^ 8);
  assign w766[55] = |(datain[91:88] ^ 11);
  assign w766[56] = |(datain[87:84] ^ 0);
  assign w766[57] = |(datain[83:80] ^ 14);
  assign w766[58] = |(datain[79:76] ^ 3);
  assign w766[59] = |(datain[75:72] ^ 10);
  assign w766[60] = |(datain[71:68] ^ 0);
  assign w766[61] = |(datain[67:64] ^ 1);
  assign w766[62] = |(datain[63:60] ^ 11);
  assign w766[63] = |(datain[59:56] ^ 10);
  assign w766[64] = |(datain[55:52] ^ 0);
  assign w766[65] = |(datain[51:48] ^ 0);
  assign w766[66] = |(datain[47:44] ^ 0);
  assign w766[67] = |(datain[43:40] ^ 5);
  assign w766[68] = |(datain[39:36] ^ 12);
  assign w766[69] = |(datain[35:32] ^ 13);
  assign w766[70] = |(datain[31:28] ^ 2);
  assign w766[71] = |(datain[27:24] ^ 1);
  assign w766[72] = |(datain[23:20] ^ 11);
  assign w766[73] = |(datain[19:16] ^ 4);
  assign w766[74] = |(datain[15:12] ^ 3);
  assign w766[75] = |(datain[11:8] ^ 14);
  assign comp[766] = ~(|w766);
  wire [62-1:0] w767;
  assign w767[0] = |(datain[311:308] ^ 6);
  assign w767[1] = |(datain[307:304] ^ 1);
  assign w767[2] = |(datain[303:300] ^ 7);
  assign w767[3] = |(datain[299:296] ^ 2);
  assign w767[4] = |(datain[295:292] ^ 6);
  assign w767[5] = |(datain[291:288] ^ 10);
  assign w767[6] = |(datain[287:284] ^ 2);
  assign w767[7] = |(datain[283:280] ^ 0);
  assign w767[8] = |(datain[279:276] ^ 6);
  assign w767[9] = |(datain[275:272] ^ 1);
  assign w767[10] = |(datain[271:268] ^ 2);
  assign w767[11] = |(datain[267:264] ^ 0);
  assign w767[12] = |(datain[263:260] ^ 2);
  assign w767[13] = |(datain[259:256] ^ 13);
  assign w767[14] = |(datain[255:252] ^ 7);
  assign w767[15] = |(datain[251:248] ^ 9);
  assign w767[16] = |(datain[247:244] ^ 2);
  assign w767[17] = |(datain[243:240] ^ 0);
  assign w767[18] = |(datain[239:236] ^ 7);
  assign w767[19] = |(datain[235:232] ^ 6);
  assign w767[20] = |(datain[231:228] ^ 5);
  assign w767[21] = |(datain[227:224] ^ 15);
  assign w767[22] = |(datain[223:220] ^ 6);
  assign w767[23] = |(datain[219:216] ^ 15);
  assign w767[24] = |(datain[215:212] ^ 5);
  assign w767[25] = |(datain[211:208] ^ 15);
  assign w767[26] = |(datain[207:204] ^ 6);
  assign w767[27] = |(datain[203:200] ^ 2);
  assign w767[28] = |(datain[199:196] ^ 6);
  assign w767[29] = |(datain[195:192] ^ 5);
  assign w767[30] = |(datain[191:188] ^ 2);
  assign w767[31] = |(datain[187:184] ^ 14);
  assign w767[32] = |(datain[183:180] ^ 6);
  assign w767[33] = |(datain[179:176] ^ 1);
  assign w767[34] = |(datain[175:172] ^ 7);
  assign w767[35] = |(datain[171:168] ^ 2);
  assign w767[36] = |(datain[167:164] ^ 6);
  assign w767[37] = |(datain[163:160] ^ 10);
  assign w767[38] = |(datain[159:156] ^ 2);
  assign w767[39] = |(datain[155:152] ^ 0);
  assign w767[40] = |(datain[151:148] ^ 7);
  assign w767[41] = |(datain[147:144] ^ 6);
  assign w767[42] = |(datain[143:140] ^ 5);
  assign w767[43] = |(datain[139:136] ^ 15);
  assign w767[44] = |(datain[135:132] ^ 6);
  assign w767[45] = |(datain[131:128] ^ 15);
  assign w767[46] = |(datain[127:124] ^ 5);
  assign w767[47] = |(datain[123:120] ^ 15);
  assign w767[48] = |(datain[119:116] ^ 6);
  assign w767[49] = |(datain[115:112] ^ 2);
  assign w767[50] = |(datain[111:108] ^ 6);
  assign w767[51] = |(datain[107:104] ^ 5);
  assign w767[52] = |(datain[103:100] ^ 2);
  assign w767[53] = |(datain[99:96] ^ 14);
  assign w767[54] = |(datain[95:92] ^ 6);
  assign w767[55] = |(datain[91:88] ^ 5);
  assign w767[56] = |(datain[87:84] ^ 7);
  assign w767[57] = |(datain[83:80] ^ 8);
  assign w767[58] = |(datain[79:76] ^ 6);
  assign w767[59] = |(datain[75:72] ^ 5);
  assign w767[60] = |(datain[71:68] ^ 2);
  assign w767[61] = |(datain[67:64] ^ 0);
  assign comp[767] = ~(|w767);
  wire [76-1:0] w768;
  assign w768[0] = |(datain[311:308] ^ 3);
  assign w768[1] = |(datain[307:304] ^ 3);
  assign w768[2] = |(datain[303:300] ^ 12);
  assign w768[3] = |(datain[299:296] ^ 0);
  assign w768[4] = |(datain[295:292] ^ 9);
  assign w768[5] = |(datain[291:288] ^ 14);
  assign w768[6] = |(datain[287:284] ^ 9);
  assign w768[7] = |(datain[283:280] ^ 15);
  assign w768[8] = |(datain[279:276] ^ 8);
  assign w768[9] = |(datain[275:272] ^ 0);
  assign w768[10] = |(datain[271:268] ^ 12);
  assign w768[11] = |(datain[267:264] ^ 4);
  assign w768[12] = |(datain[263:260] ^ 3);
  assign w768[13] = |(datain[259:256] ^ 14);
  assign w768[14] = |(datain[255:252] ^ 5);
  assign w768[15] = |(datain[251:248] ^ 0);
  assign w768[16] = |(datain[247:244] ^ 8);
  assign w768[17] = |(datain[243:240] ^ 11);
  assign w768[18] = |(datain[239:236] ^ 0);
  assign w768[19] = |(datain[235:232] ^ 14);
  assign w768[20] = |(datain[231:228] ^ 3);
  assign w768[21] = |(datain[227:224] ^ 13);
  assign w768[22] = |(datain[223:220] ^ 0);
  assign w768[23] = |(datain[219:216] ^ 1);
  assign w768[24] = |(datain[215:212] ^ 11);
  assign w768[25] = |(datain[211:208] ^ 10);
  assign w768[26] = |(datain[207:204] ^ 0);
  assign w768[27] = |(datain[203:200] ^ 0);
  assign w768[28] = |(datain[199:196] ^ 0);
  assign w768[29] = |(datain[195:192] ^ 1);
  assign w768[30] = |(datain[191:188] ^ 12);
  assign w768[31] = |(datain[187:184] ^ 13);
  assign w768[32] = |(datain[183:180] ^ 2);
  assign w768[33] = |(datain[179:176] ^ 1);
  assign w768[34] = |(datain[175:172] ^ 11);
  assign w768[35] = |(datain[171:168] ^ 8);
  assign w768[36] = |(datain[167:164] ^ 0);
  assign w768[37] = |(datain[163:160] ^ 2);
  assign w768[38] = |(datain[159:156] ^ 4);
  assign w768[39] = |(datain[155:152] ^ 2);
  assign w768[40] = |(datain[151:148] ^ 3);
  assign w768[41] = |(datain[147:144] ^ 3);
  assign w768[42] = |(datain[143:140] ^ 12);
  assign w768[43] = |(datain[139:136] ^ 9);
  assign w768[44] = |(datain[135:132] ^ 3);
  assign w768[45] = |(datain[131:128] ^ 3);
  assign w768[46] = |(datain[127:124] ^ 13);
  assign w768[47] = |(datain[123:120] ^ 2);
  assign w768[48] = |(datain[119:116] ^ 12);
  assign w768[49] = |(datain[115:112] ^ 13);
  assign w768[50] = |(datain[111:108] ^ 2);
  assign w768[51] = |(datain[107:104] ^ 1);
  assign w768[52] = |(datain[103:100] ^ 5);
  assign w768[53] = |(datain[99:96] ^ 8);
  assign w768[54] = |(datain[95:92] ^ 8);
  assign w768[55] = |(datain[91:88] ^ 11);
  assign w768[56] = |(datain[87:84] ^ 0);
  assign w768[57] = |(datain[83:80] ^ 14);
  assign w768[58] = |(datain[79:76] ^ 4);
  assign w768[59] = |(datain[75:72] ^ 1);
  assign w768[60] = |(datain[71:68] ^ 0);
  assign w768[61] = |(datain[67:64] ^ 1);
  assign w768[62] = |(datain[63:60] ^ 11);
  assign w768[63] = |(datain[59:56] ^ 10);
  assign w768[64] = |(datain[55:52] ^ 0);
  assign w768[65] = |(datain[51:48] ^ 0);
  assign w768[66] = |(datain[47:44] ^ 0);
  assign w768[67] = |(datain[43:40] ^ 5);
  assign w768[68] = |(datain[39:36] ^ 12);
  assign w768[69] = |(datain[35:32] ^ 13);
  assign w768[70] = |(datain[31:28] ^ 2);
  assign w768[71] = |(datain[27:24] ^ 1);
  assign w768[72] = |(datain[23:20] ^ 11);
  assign w768[73] = |(datain[19:16] ^ 4);
  assign w768[74] = |(datain[15:12] ^ 3);
  assign w768[75] = |(datain[11:8] ^ 14);
  assign comp[768] = ~(|w768);
  wire [72-1:0] w769;
  assign w769[0] = |(datain[311:308] ^ 2);
  assign w769[1] = |(datain[307:304] ^ 0);
  assign w769[2] = |(datain[303:300] ^ 6);
  assign w769[3] = |(datain[299:296] ^ 9);
  assign w769[4] = |(datain[295:292] ^ 6);
  assign w769[5] = |(datain[291:288] ^ 14);
  assign w769[6] = |(datain[287:284] ^ 2);
  assign w769[7] = |(datain[283:280] ^ 0);
  assign w769[8] = |(datain[279:276] ^ 2);
  assign w769[9] = |(datain[275:272] ^ 8);
  assign w769[10] = |(datain[271:268] ^ 2);
  assign w769[11] = |(datain[267:264] ^ 10);
  assign w769[12] = |(datain[263:260] ^ 2);
  assign w769[13] = |(datain[259:256] ^ 14);
  assign w769[14] = |(datain[255:252] ^ 6);
  assign w769[15] = |(datain[251:248] ^ 2);
  assign w769[16] = |(datain[247:244] ^ 6);
  assign w769[17] = |(datain[243:240] ^ 1);
  assign w769[18] = |(datain[239:236] ^ 7);
  assign w769[19] = |(datain[235:232] ^ 4);
  assign w769[20] = |(datain[231:228] ^ 2);
  assign w769[21] = |(datain[227:224] ^ 9);
  assign w769[22] = |(datain[223:220] ^ 2);
  assign w769[23] = |(datain[219:216] ^ 0);
  assign w769[24] = |(datain[215:212] ^ 6);
  assign w769[25] = |(datain[211:208] ^ 4);
  assign w769[26] = |(datain[207:204] ^ 6);
  assign w769[27] = |(datain[203:200] ^ 15);
  assign w769[28] = |(datain[199:196] ^ 2);
  assign w769[29] = |(datain[195:192] ^ 0);
  assign w769[30] = |(datain[191:188] ^ 6);
  assign w769[31] = |(datain[187:184] ^ 3);
  assign w769[32] = |(datain[183:180] ^ 6);
  assign w769[33] = |(datain[179:176] ^ 1);
  assign w769[34] = |(datain[175:172] ^ 6);
  assign w769[35] = |(datain[171:168] ^ 12);
  assign w769[36] = |(datain[167:164] ^ 6);
  assign w769[37] = |(datain[163:160] ^ 12);
  assign w769[38] = |(datain[159:156] ^ 2);
  assign w769[39] = |(datain[155:152] ^ 0);
  assign w769[40] = |(datain[151:148] ^ 2);
  assign w769[41] = |(datain[147:144] ^ 5);
  assign w769[42] = |(datain[143:140] ^ 3);
  assign w769[43] = |(datain[139:136] ^ 0);
  assign w769[44] = |(datain[135:132] ^ 2);
  assign w769[45] = |(datain[131:128] ^ 0);
  assign w769[46] = |(datain[127:124] ^ 4);
  assign w769[47] = |(datain[123:120] ^ 4);
  assign w769[48] = |(datain[119:116] ^ 6);
  assign w769[49] = |(datain[115:112] ^ 5);
  assign w769[50] = |(datain[111:108] ^ 6);
  assign w769[51] = |(datain[107:104] ^ 1);
  assign w769[52] = |(datain[103:100] ^ 6);
  assign w769[53] = |(datain[99:96] ^ 4);
  assign w769[54] = |(datain[95:92] ^ 5);
  assign w769[55] = |(datain[91:88] ^ 15);
  assign w769[56] = |(datain[87:84] ^ 4);
  assign w769[57] = |(datain[83:80] ^ 2);
  assign w769[58] = |(datain[79:76] ^ 7);
  assign w769[59] = |(datain[75:72] ^ 9);
  assign w769[60] = |(datain[71:68] ^ 7);
  assign w769[61] = |(datain[67:64] ^ 4);
  assign w769[62] = |(datain[63:60] ^ 6);
  assign w769[63] = |(datain[59:56] ^ 5);
  assign w769[64] = |(datain[55:52] ^ 2);
  assign w769[65] = |(datain[51:48] ^ 0);
  assign w769[66] = |(datain[47:44] ^ 2);
  assign w769[67] = |(datain[43:40] ^ 5);
  assign w769[68] = |(datain[39:36] ^ 2);
  assign w769[69] = |(datain[35:32] ^ 5);
  assign w769[70] = |(datain[31:28] ^ 6);
  assign w769[71] = |(datain[27:24] ^ 6);
  assign comp[769] = ~(|w769);
  wire [56-1:0] w770;
  assign w770[0] = |(datain[311:308] ^ 2);
  assign w770[1] = |(datain[307:304] ^ 14);
  assign w770[2] = |(datain[303:300] ^ 6);
  assign w770[3] = |(datain[299:296] ^ 3);
  assign w770[4] = |(datain[295:292] ^ 6);
  assign w770[5] = |(datain[291:288] ^ 15);
  assign w770[6] = |(datain[287:284] ^ 6);
  assign w770[7] = |(datain[283:280] ^ 13);
  assign w770[8] = |(datain[279:276] ^ 0);
  assign w770[9] = |(datain[275:272] ^ 13);
  assign w770[10] = |(datain[271:268] ^ 0);
  assign w770[11] = |(datain[267:264] ^ 10);
  assign w770[12] = |(datain[263:260] ^ 6);
  assign w770[13] = |(datain[259:256] ^ 4);
  assign w770[14] = |(datain[255:252] ^ 6);
  assign w770[15] = |(datain[251:248] ^ 5);
  assign w770[16] = |(datain[247:244] ^ 6);
  assign w770[17] = |(datain[243:240] ^ 12);
  assign w770[18] = |(datain[239:236] ^ 2);
  assign w770[19] = |(datain[235:232] ^ 0);
  assign w770[20] = |(datain[231:228] ^ 4);
  assign w770[21] = |(datain[227:224] ^ 3);
  assign w770[22] = |(datain[223:220] ^ 3);
  assign w770[23] = |(datain[219:216] ^ 10);
  assign w770[24] = |(datain[215:212] ^ 5);
  assign w770[25] = |(datain[211:208] ^ 12);
  assign w770[26] = |(datain[207:204] ^ 5);
  assign w770[27] = |(datain[203:200] ^ 7);
  assign w770[28] = |(datain[199:196] ^ 4);
  assign w770[29] = |(datain[195:192] ^ 9);
  assign w770[30] = |(datain[191:188] ^ 4);
  assign w770[31] = |(datain[187:184] ^ 14);
  assign w770[32] = |(datain[183:180] ^ 4);
  assign w770[33] = |(datain[179:176] ^ 4);
  assign w770[34] = |(datain[175:172] ^ 4);
  assign w770[35] = |(datain[171:168] ^ 15);
  assign w770[36] = |(datain[167:164] ^ 5);
  assign w770[37] = |(datain[163:160] ^ 7);
  assign w770[38] = |(datain[159:156] ^ 5);
  assign w770[39] = |(datain[155:152] ^ 3);
  assign w770[40] = |(datain[151:148] ^ 5);
  assign w770[41] = |(datain[147:144] ^ 12);
  assign w770[42] = |(datain[143:140] ^ 7);
  assign w770[43] = |(datain[139:136] ^ 7);
  assign w770[44] = |(datain[135:132] ^ 6);
  assign w770[45] = |(datain[131:128] ^ 9);
  assign w770[46] = |(datain[127:124] ^ 6);
  assign w770[47] = |(datain[123:120] ^ 14);
  assign w770[48] = |(datain[119:116] ^ 2);
  assign w770[49] = |(datain[115:112] ^ 14);
  assign w770[50] = |(datain[111:108] ^ 6);
  assign w770[51] = |(datain[107:104] ^ 3);
  assign w770[52] = |(datain[103:100] ^ 6);
  assign w770[53] = |(datain[99:96] ^ 15);
  assign w770[54] = |(datain[95:92] ^ 6);
  assign w770[55] = |(datain[91:88] ^ 13);
  assign comp[770] = ~(|w770);
  wire [44-1:0] w771;
  assign w771[0] = |(datain[311:308] ^ 6);
  assign w771[1] = |(datain[307:304] ^ 5);
  assign w771[2] = |(datain[303:300] ^ 6);
  assign w771[3] = |(datain[299:296] ^ 3);
  assign w771[4] = |(datain[295:292] ^ 6);
  assign w771[5] = |(datain[291:288] ^ 8);
  assign w771[6] = |(datain[287:284] ^ 6);
  assign w771[7] = |(datain[283:280] ^ 15);
  assign w771[8] = |(datain[279:276] ^ 2);
  assign w771[9] = |(datain[275:272] ^ 0);
  assign w771[10] = |(datain[271:268] ^ 2);
  assign w771[11] = |(datain[267:264] ^ 14);
  assign w771[12] = |(datain[263:260] ^ 4);
  assign w771[13] = |(datain[259:256] ^ 2);
  assign w771[14] = |(datain[255:252] ^ 4);
  assign w771[15] = |(datain[251:248] ^ 1);
  assign w771[16] = |(datain[247:244] ^ 5);
  assign w771[17] = |(datain[243:240] ^ 4);
  assign w771[18] = |(datain[239:236] ^ 2);
  assign w771[19] = |(datain[235:232] ^ 0);
  assign w771[20] = |(datain[231:228] ^ 7);
  assign w771[21] = |(datain[227:224] ^ 6);
  assign w771[22] = |(datain[223:220] ^ 6);
  assign w771[23] = |(datain[219:216] ^ 9);
  assign w771[24] = |(datain[215:212] ^ 7);
  assign w771[25] = |(datain[211:208] ^ 2);
  assign w771[26] = |(datain[207:204] ^ 7);
  assign w771[27] = |(datain[203:200] ^ 5);
  assign w771[28] = |(datain[199:196] ^ 7);
  assign w771[29] = |(datain[195:192] ^ 3);
  assign w771[30] = |(datain[191:188] ^ 2);
  assign w771[31] = |(datain[187:184] ^ 0);
  assign w771[32] = |(datain[183:180] ^ 2);
  assign w771[33] = |(datain[179:176] ^ 7);
  assign w771[34] = |(datain[175:172] ^ 4);
  assign w771[35] = |(datain[171:168] ^ 0);
  assign w771[36] = |(datain[167:164] ^ 4);
  assign w771[37] = |(datain[163:160] ^ 0);
  assign w771[38] = |(datain[159:156] ^ 2);
  assign w771[39] = |(datain[155:152] ^ 7);
  assign w771[40] = |(datain[151:148] ^ 2);
  assign w771[41] = |(datain[147:144] ^ 0);
  assign w771[42] = |(datain[143:140] ^ 7);
  assign w771[43] = |(datain[139:136] ^ 6);
  assign comp[771] = ~(|w771);
  wire [62-1:0] w772;
  assign w772[0] = |(datain[311:308] ^ 7);
  assign w772[1] = |(datain[307:304] ^ 10);
  assign w772[2] = |(datain[303:300] ^ 2);
  assign w772[3] = |(datain[299:296] ^ 0);
  assign w772[4] = |(datain[295:292] ^ 5);
  assign w772[5] = |(datain[291:288] ^ 11);
  assign w772[6] = |(datain[287:284] ^ 4);
  assign w772[7] = |(datain[283:280] ^ 1);
  assign w772[8] = |(datain[279:276] ^ 4);
  assign w772[9] = |(datain[275:272] ^ 2);
  assign w772[10] = |(datain[271:268] ^ 4);
  assign w772[11] = |(datain[267:264] ^ 13);
  assign w772[12] = |(datain[263:260] ^ 2);
  assign w772[13] = |(datain[259:256] ^ 0);
  assign w772[14] = |(datain[255:252] ^ 3);
  assign w772[15] = |(datain[251:248] ^ 1);
  assign w772[16] = |(datain[247:244] ^ 2);
  assign w772[17] = |(datain[243:240] ^ 14);
  assign w772[18] = |(datain[239:236] ^ 3);
  assign w772[19] = |(datain[235:232] ^ 3);
  assign w772[20] = |(datain[231:228] ^ 2);
  assign w772[21] = |(datain[227:224] ^ 0);
  assign w772[22] = |(datain[223:220] ^ 6);
  assign w772[23] = |(datain[219:216] ^ 4);
  assign w772[24] = |(datain[215:212] ^ 6);
  assign w772[25] = |(datain[211:208] ^ 5);
  assign w772[26] = |(datain[207:204] ^ 6);
  assign w772[27] = |(datain[203:200] ^ 13);
  assign w772[28] = |(datain[199:196] ^ 6);
  assign w772[29] = |(datain[195:192] ^ 15);
  assign w772[30] = |(datain[191:188] ^ 5);
  assign w772[31] = |(datain[187:184] ^ 13);
  assign w772[32] = |(datain[183:180] ^ 2);
  assign w772[33] = |(datain[179:176] ^ 0);
  assign w772[34] = |(datain[175:172] ^ 6);
  assign w772[35] = |(datain[171:168] ^ 2);
  assign w772[36] = |(datain[167:164] ^ 7);
  assign w772[37] = |(datain[163:160] ^ 9);
  assign w772[38] = |(datain[159:156] ^ 2);
  assign w772[39] = |(datain[155:152] ^ 0);
  assign w772[40] = |(datain[151:148] ^ 4);
  assign w772[41] = |(datain[147:144] ^ 4);
  assign w772[42] = |(datain[143:140] ^ 7);
  assign w772[43] = |(datain[139:136] ^ 5);
  assign w772[44] = |(datain[135:132] ^ 6);
  assign w772[45] = |(datain[131:128] ^ 11);
  assign w772[46] = |(datain[127:124] ^ 6);
  assign w772[47] = |(datain[123:120] ^ 5);
  assign w772[48] = |(datain[119:116] ^ 2);
  assign w772[49] = |(datain[115:112] ^ 15);
  assign w772[50] = |(datain[111:108] ^ 5);
  assign w772[51] = |(datain[107:104] ^ 3);
  assign w772[52] = |(datain[103:100] ^ 4);
  assign w772[53] = |(datain[99:96] ^ 13);
  assign w772[54] = |(datain[95:92] ^ 4);
  assign w772[55] = |(datain[91:88] ^ 6);
  assign w772[56] = |(datain[87:84] ^ 2);
  assign w772[57] = |(datain[83:80] ^ 5);
  assign w772[58] = |(datain[79:76] ^ 2);
  assign w772[59] = |(datain[75:72] ^ 5);
  assign w772[60] = |(datain[71:68] ^ 0);
  assign w772[61] = |(datain[67:64] ^ 13);
  assign comp[772] = ~(|w772);
  wire [76-1:0] w773;
  assign w773[0] = |(datain[311:308] ^ 2);
  assign w773[1] = |(datain[307:304] ^ 5);
  assign w773[2] = |(datain[303:300] ^ 4);
  assign w773[3] = |(datain[299:296] ^ 4);
  assign w773[4] = |(datain[295:292] ^ 7);
  assign w773[5] = |(datain[291:288] ^ 5);
  assign w773[6] = |(datain[287:284] ^ 6);
  assign w773[7] = |(datain[283:280] ^ 11);
  assign w773[8] = |(datain[279:276] ^ 6);
  assign w773[9] = |(datain[275:272] ^ 5);
  assign w773[10] = |(datain[271:268] ^ 6);
  assign w773[11] = |(datain[267:264] ^ 6);
  assign w773[12] = |(datain[263:260] ^ 2);
  assign w773[13] = |(datain[259:256] ^ 5);
  assign w773[14] = |(datain[255:252] ^ 7);
  assign w773[15] = |(datain[251:248] ^ 3);
  assign w773[16] = |(datain[247:244] ^ 6);
  assign w773[17] = |(datain[243:240] ^ 5);
  assign w773[18] = |(datain[239:236] ^ 7);
  assign w773[19] = |(datain[235:232] ^ 4);
  assign w773[20] = |(datain[231:228] ^ 2);
  assign w773[21] = |(datain[227:224] ^ 0);
  assign w773[22] = |(datain[223:220] ^ 7);
  assign w773[23] = |(datain[219:216] ^ 9);
  assign w773[24] = |(datain[215:212] ^ 6);
  assign w773[25] = |(datain[211:208] ^ 3);
  assign w773[26] = |(datain[207:204] ^ 3);
  assign w773[27] = |(datain[203:200] ^ 13);
  assign w773[28] = |(datain[199:196] ^ 6);
  assign w773[29] = |(datain[195:192] ^ 14);
  assign w773[30] = |(datain[191:188] ^ 7);
  assign w773[31] = |(datain[187:184] ^ 5);
  assign w773[32] = |(datain[183:180] ^ 6);
  assign w773[33] = |(datain[179:176] ^ 12);
  assign w773[34] = |(datain[175:172] ^ 0);
  assign w773[35] = |(datain[171:168] ^ 13);
  assign w773[36] = |(datain[167:164] ^ 0);
  assign w773[37] = |(datain[163:160] ^ 10);
  assign w773[38] = |(datain[159:156] ^ 7);
  assign w773[39] = |(datain[155:152] ^ 3);
  assign w773[40] = |(datain[151:148] ^ 6);
  assign w773[41] = |(datain[147:144] ^ 5);
  assign w773[42] = |(datain[143:140] ^ 7);
  assign w773[43] = |(datain[139:136] ^ 4);
  assign w773[44] = |(datain[135:132] ^ 2);
  assign w773[45] = |(datain[131:128] ^ 0);
  assign w773[46] = |(datain[127:124] ^ 7);
  assign w773[47] = |(datain[123:120] ^ 9);
  assign w773[48] = |(datain[119:116] ^ 6);
  assign w773[49] = |(datain[115:112] ^ 3);
  assign w773[50] = |(datain[111:108] ^ 2);
  assign w773[51] = |(datain[107:104] ^ 5);
  assign w773[52] = |(datain[103:100] ^ 4);
  assign w773[53] = |(datain[99:96] ^ 4);
  assign w773[54] = |(datain[95:92] ^ 7);
  assign w773[55] = |(datain[91:88] ^ 5);
  assign w773[56] = |(datain[87:84] ^ 6);
  assign w773[57] = |(datain[83:80] ^ 11);
  assign w773[58] = |(datain[79:76] ^ 6);
  assign w773[59] = |(datain[75:72] ^ 5);
  assign w773[60] = |(datain[71:68] ^ 6);
  assign w773[61] = |(datain[67:64] ^ 11);
  assign w773[62] = |(datain[63:60] ^ 2);
  assign w773[63] = |(datain[59:56] ^ 5);
  assign w773[64] = |(datain[55:52] ^ 3);
  assign w773[65] = |(datain[51:48] ^ 13);
  assign w773[66] = |(datain[47:44] ^ 2);
  assign w773[67] = |(datain[43:40] ^ 5);
  assign w773[68] = |(datain[39:36] ^ 7);
  assign w773[69] = |(datain[35:32] ^ 9);
  assign w773[70] = |(datain[31:28] ^ 6);
  assign w773[71] = |(datain[27:24] ^ 3);
  assign w773[72] = |(datain[23:20] ^ 2);
  assign w773[73] = |(datain[19:16] ^ 5);
  assign w773[74] = |(datain[15:12] ^ 0);
  assign w773[75] = |(datain[11:8] ^ 13);
  assign comp[773] = ~(|w773);
  wire [56-1:0] w774;
  assign w774[0] = |(datain[311:308] ^ 2);
  assign w774[1] = |(datain[307:304] ^ 10);
  assign w774[2] = |(datain[303:300] ^ 2);
  assign w774[3] = |(datain[299:296] ^ 14);
  assign w774[4] = |(datain[295:292] ^ 6);
  assign w774[5] = |(datain[291:288] ^ 2);
  assign w774[6] = |(datain[287:284] ^ 6);
  assign w774[7] = |(datain[283:280] ^ 1);
  assign w774[8] = |(datain[279:276] ^ 7);
  assign w774[9] = |(datain[275:272] ^ 4);
  assign w774[10] = |(datain[271:268] ^ 2);
  assign w774[11] = |(datain[267:264] ^ 9);
  assign w774[12] = |(datain[263:260] ^ 2);
  assign w774[13] = |(datain[259:256] ^ 0);
  assign w774[14] = |(datain[255:252] ^ 6);
  assign w774[15] = |(datain[251:248] ^ 4);
  assign w774[16] = |(datain[247:244] ^ 6);
  assign w774[17] = |(datain[243:240] ^ 15);
  assign w774[18] = |(datain[239:236] ^ 2);
  assign w774[19] = |(datain[235:232] ^ 0);
  assign w774[20] = |(datain[231:228] ^ 6);
  assign w774[21] = |(datain[227:224] ^ 3);
  assign w774[22] = |(datain[223:220] ^ 6);
  assign w774[23] = |(datain[219:216] ^ 1);
  assign w774[24] = |(datain[215:212] ^ 6);
  assign w774[25] = |(datain[211:208] ^ 12);
  assign w774[26] = |(datain[207:204] ^ 6);
  assign w774[27] = |(datain[203:200] ^ 12);
  assign w774[28] = |(datain[199:196] ^ 2);
  assign w774[29] = |(datain[195:192] ^ 0);
  assign w774[30] = |(datain[191:188] ^ 2);
  assign w774[31] = |(datain[187:184] ^ 5);
  assign w774[32] = |(datain[183:180] ^ 3);
  assign w774[33] = |(datain[179:176] ^ 0);
  assign w774[34] = |(datain[175:172] ^ 2);
  assign w774[35] = |(datain[171:168] ^ 0);
  assign w774[36] = |(datain[167:164] ^ 2);
  assign w774[37] = |(datain[163:160] ^ 15);
  assign w774[38] = |(datain[159:156] ^ 6);
  assign w774[39] = |(datain[155:152] ^ 8);
  assign w774[40] = |(datain[151:148] ^ 6);
  assign w774[41] = |(datain[147:144] ^ 1);
  assign w774[42] = |(datain[143:140] ^ 6);
  assign w774[43] = |(datain[139:136] ^ 10);
  assign w774[44] = |(datain[135:132] ^ 5);
  assign w774[45] = |(datain[131:128] ^ 15);
  assign w774[46] = |(datain[127:124] ^ 7);
  assign w774[47] = |(datain[123:120] ^ 0);
  assign w774[48] = |(datain[119:116] ^ 2);
  assign w774[49] = |(datain[115:112] ^ 0);
  assign w774[50] = |(datain[111:108] ^ 2);
  assign w774[51] = |(datain[107:104] ^ 5);
  assign w774[52] = |(datain[103:100] ^ 2);
  assign w774[53] = |(datain[99:96] ^ 5);
  assign w774[54] = |(datain[95:92] ^ 6);
  assign w774[55] = |(datain[91:88] ^ 1);
  assign comp[774] = ~(|w774);
  wire [74-1:0] w775;
  assign w775[0] = |(datain[311:308] ^ 6);
  assign w775[1] = |(datain[307:304] ^ 6);
  assign w775[2] = |(datain[303:300] ^ 6);
  assign w775[3] = |(datain[299:296] ^ 15);
  assign w775[4] = |(datain[295:292] ^ 7);
  assign w775[5] = |(datain[291:288] ^ 2);
  assign w775[6] = |(datain[287:284] ^ 2);
  assign w775[7] = |(datain[283:280] ^ 0);
  assign w775[8] = |(datain[279:276] ^ 2);
  assign w775[9] = |(datain[275:272] ^ 5);
  assign w775[10] = |(datain[271:268] ^ 2);
  assign w775[11] = |(datain[267:264] ^ 5);
  assign w775[12] = |(datain[263:260] ^ 6);
  assign w775[13] = |(datain[259:256] ^ 6);
  assign w775[14] = |(datain[255:252] ^ 2);
  assign w775[15] = |(datain[251:248] ^ 0);
  assign w775[16] = |(datain[247:244] ^ 6);
  assign w775[17] = |(datain[243:240] ^ 9);
  assign w775[18] = |(datain[239:236] ^ 6);
  assign w775[19] = |(datain[235:232] ^ 14);
  assign w775[20] = |(datain[231:228] ^ 2);
  assign w775[21] = |(datain[227:224] ^ 0);
  assign w775[22] = |(datain[223:220] ^ 2);
  assign w775[23] = |(datain[219:216] ^ 8);
  assign w775[24] = |(datain[215:212] ^ 2);
  assign w775[25] = |(datain[211:208] ^ 10);
  assign w775[26] = |(datain[207:204] ^ 2);
  assign w775[27] = |(datain[203:200] ^ 14);
  assign w775[28] = |(datain[199:196] ^ 6);
  assign w775[29] = |(datain[195:192] ^ 5);
  assign w775[30] = |(datain[191:188] ^ 7);
  assign w775[31] = |(datain[187:184] ^ 8);
  assign w775[32] = |(datain[183:180] ^ 6);
  assign w775[33] = |(datain[179:176] ^ 5);
  assign w775[34] = |(datain[175:172] ^ 2);
  assign w775[35] = |(datain[171:168] ^ 0);
  assign w775[36] = |(datain[167:164] ^ 2);
  assign w775[37] = |(datain[163:160] ^ 10);
  assign w775[38] = |(datain[159:156] ^ 2);
  assign w775[39] = |(datain[155:152] ^ 14);
  assign w775[40] = |(datain[151:148] ^ 6);
  assign w775[41] = |(datain[147:144] ^ 3);
  assign w775[42] = |(datain[143:140] ^ 6);
  assign w775[43] = |(datain[139:136] ^ 15);
  assign w775[44] = |(datain[135:132] ^ 6);
  assign w775[45] = |(datain[131:128] ^ 13);
  assign w775[46] = |(datain[127:124] ^ 2);
  assign w775[47] = |(datain[123:120] ^ 9);
  assign w775[48] = |(datain[119:116] ^ 2);
  assign w775[49] = |(datain[115:112] ^ 0);
  assign w775[50] = |(datain[111:108] ^ 6);
  assign w775[51] = |(datain[107:104] ^ 4);
  assign w775[52] = |(datain[103:100] ^ 6);
  assign w775[53] = |(datain[99:96] ^ 15);
  assign w775[54] = |(datain[95:92] ^ 2);
  assign w775[55] = |(datain[91:88] ^ 0);
  assign w775[56] = |(datain[87:84] ^ 7);
  assign w775[57] = |(datain[83:80] ^ 3);
  assign w775[58] = |(datain[79:76] ^ 6);
  assign w775[59] = |(datain[75:72] ^ 5);
  assign w775[60] = |(datain[71:68] ^ 7);
  assign w775[61] = |(datain[67:64] ^ 4);
  assign w775[62] = |(datain[63:60] ^ 2);
  assign w775[63] = |(datain[59:56] ^ 0);
  assign w775[64] = |(datain[55:52] ^ 4);
  assign w775[65] = |(datain[51:48] ^ 1);
  assign w775[66] = |(datain[47:44] ^ 3);
  assign w775[67] = |(datain[43:40] ^ 13);
  assign w775[68] = |(datain[39:36] ^ 2);
  assign w775[69] = |(datain[35:32] ^ 5);
  assign w775[70] = |(datain[31:28] ^ 2);
  assign w775[71] = |(datain[27:24] ^ 5);
  assign w775[72] = |(datain[23:20] ^ 6);
  assign w775[73] = |(datain[19:16] ^ 6);
  assign comp[775] = ~(|w775);
  wire [76-1:0] w776;
  assign w776[0] = |(datain[311:308] ^ 3);
  assign w776[1] = |(datain[307:304] ^ 15);
  assign w776[2] = |(datain[303:300] ^ 2);
  assign w776[3] = |(datain[299:296] ^ 14);
  assign w776[4] = |(datain[295:292] ^ 8);
  assign w776[5] = |(datain[291:288] ^ 11);
  assign w776[6] = |(datain[287:284] ^ 1);
  assign w776[7] = |(datain[283:280] ^ 14);
  assign w776[8] = |(datain[279:276] ^ 1);
  assign w776[9] = |(datain[275:272] ^ 2);
  assign w776[10] = |(datain[271:268] ^ 0);
  assign w776[11] = |(datain[267:264] ^ 1);
  assign w776[12] = |(datain[263:260] ^ 12);
  assign w776[13] = |(datain[259:256] ^ 13);
  assign w776[14] = |(datain[255:252] ^ 15);
  assign w776[15] = |(datain[251:248] ^ 1);
  assign w776[16] = |(datain[247:244] ^ 12);
  assign w776[17] = |(datain[243:240] ^ 3);
  assign w776[18] = |(datain[239:236] ^ 11);
  assign w776[19] = |(datain[235:232] ^ 4);
  assign w776[20] = |(datain[231:228] ^ 4);
  assign w776[21] = |(datain[227:224] ^ 0);
  assign w776[22] = |(datain[223:220] ^ 2);
  assign w776[23] = |(datain[219:216] ^ 14);
  assign w776[24] = |(datain[215:212] ^ 8);
  assign w776[25] = |(datain[211:208] ^ 11);
  assign w776[26] = |(datain[207:204] ^ 1);
  assign w776[27] = |(datain[203:200] ^ 14);
  assign w776[28] = |(datain[199:196] ^ 1);
  assign w776[29] = |(datain[195:192] ^ 2);
  assign w776[30] = |(datain[191:188] ^ 0);
  assign w776[31] = |(datain[187:184] ^ 1);
  assign w776[32] = |(datain[183:180] ^ 12);
  assign w776[33] = |(datain[179:176] ^ 13);
  assign w776[34] = |(datain[175:172] ^ 15);
  assign w776[35] = |(datain[171:168] ^ 1);
  assign w776[36] = |(datain[167:164] ^ 12);
  assign w776[37] = |(datain[163:160] ^ 3);
  assign w776[38] = |(datain[159:156] ^ 11);
  assign w776[39] = |(datain[155:152] ^ 0);
  assign w776[40] = |(datain[151:148] ^ 0);
  assign w776[41] = |(datain[147:144] ^ 0);
  assign w776[42] = |(datain[143:140] ^ 12);
  assign w776[43] = |(datain[139:136] ^ 15);
  assign w776[44] = |(datain[135:132] ^ 2);
  assign w776[45] = |(datain[131:128] ^ 14);
  assign w776[46] = |(datain[127:124] ^ 8);
  assign w776[47] = |(datain[123:120] ^ 0);
  assign w776[48] = |(datain[119:116] ^ 3);
  assign w776[49] = |(datain[115:112] ^ 14);
  assign w776[50] = |(datain[111:108] ^ 4);
  assign w776[51] = |(datain[107:104] ^ 15);
  assign w776[52] = |(datain[103:100] ^ 0);
  assign w776[53] = |(datain[99:96] ^ 1);
  assign w776[54] = |(datain[95:92] ^ 2);
  assign w776[55] = |(datain[91:88] ^ 0);
  assign w776[56] = |(datain[87:84] ^ 7);
  assign w776[57] = |(datain[83:80] ^ 5);
  assign w776[58] = |(datain[79:76] ^ 0);
  assign w776[59] = |(datain[75:72] ^ 9);
  assign w776[60] = |(datain[71:68] ^ 14);
  assign w776[61] = |(datain[67:64] ^ 8);
  assign w776[62] = |(datain[63:60] ^ 6);
  assign w776[63] = |(datain[59:56] ^ 1);
  assign w776[64] = |(datain[55:52] ^ 0);
  assign w776[65] = |(datain[51:48] ^ 1);
  assign w776[66] = |(datain[47:44] ^ 2);
  assign w776[67] = |(datain[43:40] ^ 14);
  assign w776[68] = |(datain[39:36] ^ 12);
  assign w776[69] = |(datain[35:32] ^ 6);
  assign w776[70] = |(datain[31:28] ^ 0);
  assign w776[71] = |(datain[27:24] ^ 6);
  assign w776[72] = |(datain[23:20] ^ 4);
  assign w776[73] = |(datain[19:16] ^ 15);
  assign w776[74] = |(datain[15:12] ^ 0);
  assign w776[75] = |(datain[11:8] ^ 1);
  assign comp[776] = ~(|w776);
  wire [72-1:0] w777;
  assign w777[0] = |(datain[311:308] ^ 2);
  assign w777[1] = |(datain[307:304] ^ 0);
  assign w777[2] = |(datain[303:300] ^ 6);
  assign w777[3] = |(datain[299:296] ^ 9);
  assign w777[4] = |(datain[295:292] ^ 6);
  assign w777[5] = |(datain[291:288] ^ 14);
  assign w777[6] = |(datain[287:284] ^ 2);
  assign w777[7] = |(datain[283:280] ^ 0);
  assign w777[8] = |(datain[279:276] ^ 2);
  assign w777[9] = |(datain[275:272] ^ 8);
  assign w777[10] = |(datain[271:268] ^ 2);
  assign w777[11] = |(datain[267:264] ^ 10);
  assign w777[12] = |(datain[263:260] ^ 2);
  assign w777[13] = |(datain[259:256] ^ 14);
  assign w777[14] = |(datain[255:252] ^ 6);
  assign w777[15] = |(datain[251:248] ^ 2);
  assign w777[16] = |(datain[247:244] ^ 6);
  assign w777[17] = |(datain[243:240] ^ 1);
  assign w777[18] = |(datain[239:236] ^ 7);
  assign w777[19] = |(datain[235:232] ^ 4);
  assign w777[20] = |(datain[231:228] ^ 2);
  assign w777[21] = |(datain[227:224] ^ 9);
  assign w777[22] = |(datain[223:220] ^ 2);
  assign w777[23] = |(datain[219:216] ^ 0);
  assign w777[24] = |(datain[215:212] ^ 6);
  assign w777[25] = |(datain[211:208] ^ 4);
  assign w777[26] = |(datain[207:204] ^ 6);
  assign w777[27] = |(datain[203:200] ^ 15);
  assign w777[28] = |(datain[199:196] ^ 2);
  assign w777[29] = |(datain[195:192] ^ 0);
  assign w777[30] = |(datain[191:188] ^ 6);
  assign w777[31] = |(datain[187:184] ^ 3);
  assign w777[32] = |(datain[183:180] ^ 6);
  assign w777[33] = |(datain[179:176] ^ 1);
  assign w777[34] = |(datain[175:172] ^ 6);
  assign w777[35] = |(datain[171:168] ^ 12);
  assign w777[36] = |(datain[167:164] ^ 6);
  assign w777[37] = |(datain[163:160] ^ 12);
  assign w777[38] = |(datain[159:156] ^ 2);
  assign w777[39] = |(datain[155:152] ^ 0);
  assign w777[40] = |(datain[151:148] ^ 2);
  assign w777[41] = |(datain[147:144] ^ 5);
  assign w777[42] = |(datain[143:140] ^ 3);
  assign w777[43] = |(datain[139:136] ^ 0);
  assign w777[44] = |(datain[135:132] ^ 2);
  assign w777[45] = |(datain[131:128] ^ 0);
  assign w777[46] = |(datain[127:124] ^ 5);
  assign w777[47] = |(datain[123:120] ^ 0);
  assign w777[48] = |(datain[119:116] ^ 5);
  assign w777[49] = |(datain[115:112] ^ 5);
  assign w777[50] = |(datain[111:108] ^ 5);
  assign w777[51] = |(datain[107:104] ^ 3);
  assign w777[52] = |(datain[103:100] ^ 4);
  assign w777[53] = |(datain[99:96] ^ 8);
  assign w777[54] = |(datain[95:92] ^ 4);
  assign w777[55] = |(datain[91:88] ^ 9);
  assign w777[56] = |(datain[87:84] ^ 5);
  assign w777[57] = |(datain[83:80] ^ 3);
  assign w777[58] = |(datain[79:76] ^ 5);
  assign w777[59] = |(datain[75:72] ^ 4);
  assign w777[60] = |(datain[71:68] ^ 4);
  assign w777[61] = |(datain[67:64] ^ 9);
  assign w777[62] = |(datain[63:60] ^ 4);
  assign w777[63] = |(datain[59:56] ^ 11);
  assign w777[64] = |(datain[55:52] ^ 2);
  assign w777[65] = |(datain[51:48] ^ 0);
  assign w777[66] = |(datain[47:44] ^ 2);
  assign w777[67] = |(datain[43:40] ^ 5);
  assign w777[68] = |(datain[39:36] ^ 2);
  assign w777[69] = |(datain[35:32] ^ 5);
  assign w777[70] = |(datain[31:28] ^ 6);
  assign w777[71] = |(datain[27:24] ^ 6);
  assign comp[777] = ~(|w777);
  wire [34-1:0] w778;
  assign w778[0] = |(datain[311:308] ^ 5);
  assign w778[1] = |(datain[307:304] ^ 7);
  assign w778[2] = |(datain[303:300] ^ 11);
  assign w778[3] = |(datain[299:296] ^ 4);
  assign w778[4] = |(datain[295:292] ^ 0);
  assign w778[5] = |(datain[291:288] ^ 11);
  assign w778[6] = |(datain[287:284] ^ 12);
  assign w778[7] = |(datain[283:280] ^ 13);
  assign w778[8] = |(datain[279:276] ^ 2);
  assign w778[9] = |(datain[275:272] ^ 1);
  assign w778[10] = |(datain[271:268] ^ 0);
  assign w778[11] = |(datain[267:264] ^ 10);
  assign w778[12] = |(datain[263:260] ^ 12);
  assign w778[13] = |(datain[259:256] ^ 0);
  assign w778[14] = |(datain[255:252] ^ 7);
  assign w778[15] = |(datain[251:248] ^ 5);
  assign w778[16] = |(datain[247:244] ^ 0);
  assign w778[17] = |(datain[243:240] ^ 2);
  assign w778[18] = |(datain[239:236] ^ 12);
  assign w778[19] = |(datain[235:232] ^ 13);
  assign w778[20] = |(datain[231:228] ^ 2);
  assign w778[21] = |(datain[227:224] ^ 0);
  assign w778[22] = |(datain[223:220] ^ 11);
  assign w778[23] = |(datain[219:216] ^ 4);
  assign w778[24] = |(datain[215:212] ^ 0);
  assign w778[25] = |(datain[211:208] ^ 6);
  assign w778[26] = |(datain[207:204] ^ 11);
  assign w778[27] = |(datain[203:200] ^ 2);
  assign w778[28] = |(datain[199:196] ^ 15);
  assign w778[29] = |(datain[195:192] ^ 15);
  assign w778[30] = |(datain[191:188] ^ 12);
  assign w778[31] = |(datain[187:184] ^ 13);
  assign w778[32] = |(datain[183:180] ^ 2);
  assign w778[33] = |(datain[179:176] ^ 1);
  assign comp[778] = ~(|w778);
  wire [60-1:0] w779;
  assign w779[0] = |(datain[311:308] ^ 7);
  assign w779[1] = |(datain[307:304] ^ 2);
  assign w779[2] = |(datain[303:300] ^ 2);
  assign w779[3] = |(datain[299:296] ^ 0);
  assign w779[4] = |(datain[295:292] ^ 2);
  assign w779[5] = |(datain[291:288] ^ 5);
  assign w779[6] = |(datain[287:284] ^ 2);
  assign w779[7] = |(datain[283:280] ^ 5);
  assign w779[8] = |(datain[279:276] ^ 6);
  assign w779[9] = |(datain[275:272] ^ 2);
  assign w779[10] = |(datain[271:268] ^ 2);
  assign w779[11] = |(datain[267:264] ^ 0);
  assign w779[12] = |(datain[263:260] ^ 6);
  assign w779[13] = |(datain[259:256] ^ 9);
  assign w779[14] = |(datain[255:252] ^ 6);
  assign w779[15] = |(datain[251:248] ^ 14);
  assign w779[16] = |(datain[247:244] ^ 2);
  assign w779[17] = |(datain[243:240] ^ 0);
  assign w779[18] = |(datain[239:236] ^ 2);
  assign w779[19] = |(datain[235:232] ^ 8);
  assign w779[20] = |(datain[231:228] ^ 2);
  assign w779[21] = |(datain[227:224] ^ 10);
  assign w779[22] = |(datain[223:220] ^ 2);
  assign w779[23] = |(datain[219:216] ^ 14);
  assign w779[24] = |(datain[215:212] ^ 6);
  assign w779[25] = |(datain[211:208] ^ 2);
  assign w779[26] = |(datain[207:204] ^ 2);
  assign w779[27] = |(datain[203:200] ^ 10);
  assign w779[28] = |(datain[199:196] ^ 2);
  assign w779[29] = |(datain[195:192] ^ 9);
  assign w779[30] = |(datain[191:188] ^ 2);
  assign w779[31] = |(datain[187:184] ^ 0);
  assign w779[32] = |(datain[183:180] ^ 6);
  assign w779[33] = |(datain[179:176] ^ 4);
  assign w779[34] = |(datain[175:172] ^ 6);
  assign w779[35] = |(datain[171:168] ^ 15);
  assign w779[36] = |(datain[167:164] ^ 2);
  assign w779[37] = |(datain[163:160] ^ 0);
  assign w779[38] = |(datain[159:156] ^ 6);
  assign w779[39] = |(datain[155:152] ^ 3);
  assign w779[40] = |(datain[151:148] ^ 6);
  assign w779[41] = |(datain[147:144] ^ 15);
  assign w779[42] = |(datain[143:140] ^ 7);
  assign w779[43] = |(datain[139:136] ^ 0);
  assign w779[44] = |(datain[135:132] ^ 7);
  assign w779[45] = |(datain[131:128] ^ 9);
  assign w779[46] = |(datain[127:124] ^ 2);
  assign w779[47] = |(datain[123:120] ^ 0);
  assign w779[48] = |(datain[119:116] ^ 2);
  assign w779[49] = |(datain[115:112] ^ 5);
  assign w779[50] = |(datain[111:108] ^ 3);
  assign w779[51] = |(datain[107:104] ^ 0);
  assign w779[52] = |(datain[103:100] ^ 2);
  assign w779[53] = |(datain[99:96] ^ 0);
  assign w779[54] = |(datain[95:92] ^ 2);
  assign w779[55] = |(datain[91:88] ^ 5);
  assign w779[56] = |(datain[87:84] ^ 2);
  assign w779[57] = |(datain[83:80] ^ 5);
  assign w779[58] = |(datain[79:76] ^ 6);
  assign w779[59] = |(datain[75:72] ^ 2);
  assign comp[779] = ~(|w779);
  wire [62-1:0] w780;
  assign w780[0] = |(datain[311:308] ^ 6);
  assign w780[1] = |(datain[307:304] ^ 15);
  assign w780[2] = |(datain[303:300] ^ 7);
  assign w780[3] = |(datain[299:296] ^ 2);
  assign w780[4] = |(datain[295:292] ^ 2);
  assign w780[5] = |(datain[291:288] ^ 0);
  assign w780[6] = |(datain[287:284] ^ 2);
  assign w780[7] = |(datain[283:280] ^ 5);
  assign w780[8] = |(datain[279:276] ^ 2);
  assign w780[9] = |(datain[275:272] ^ 5);
  assign w780[10] = |(datain[271:268] ^ 6);
  assign w780[11] = |(datain[267:264] ^ 2);
  assign w780[12] = |(datain[263:260] ^ 2);
  assign w780[13] = |(datain[259:256] ^ 0);
  assign w780[14] = |(datain[255:252] ^ 6);
  assign w780[15] = |(datain[251:248] ^ 9);
  assign w780[16] = |(datain[247:244] ^ 6);
  assign w780[17] = |(datain[243:240] ^ 14);
  assign w780[18] = |(datain[239:236] ^ 2);
  assign w780[19] = |(datain[235:232] ^ 0);
  assign w780[20] = |(datain[231:228] ^ 2);
  assign w780[21] = |(datain[227:224] ^ 8);
  assign w780[22] = |(datain[223:220] ^ 2);
  assign w780[23] = |(datain[219:216] ^ 10);
  assign w780[24] = |(datain[215:212] ^ 2);
  assign w780[25] = |(datain[211:208] ^ 14);
  assign w780[26] = |(datain[207:204] ^ 6);
  assign w780[27] = |(datain[203:200] ^ 2);
  assign w780[28] = |(datain[199:196] ^ 2);
  assign w780[29] = |(datain[195:192] ^ 10);
  assign w780[30] = |(datain[191:188] ^ 2);
  assign w780[31] = |(datain[187:184] ^ 9);
  assign w780[32] = |(datain[183:180] ^ 2);
  assign w780[33] = |(datain[179:176] ^ 0);
  assign w780[34] = |(datain[175:172] ^ 6);
  assign w780[35] = |(datain[171:168] ^ 4);
  assign w780[36] = |(datain[167:164] ^ 6);
  assign w780[37] = |(datain[163:160] ^ 15);
  assign w780[38] = |(datain[159:156] ^ 2);
  assign w780[39] = |(datain[155:152] ^ 0);
  assign w780[40] = |(datain[151:148] ^ 6);
  assign w780[41] = |(datain[147:144] ^ 3);
  assign w780[42] = |(datain[143:140] ^ 6);
  assign w780[43] = |(datain[139:136] ^ 15);
  assign w780[44] = |(datain[135:132] ^ 7);
  assign w780[45] = |(datain[131:128] ^ 0);
  assign w780[46] = |(datain[127:124] ^ 7);
  assign w780[47] = |(datain[123:120] ^ 9);
  assign w780[48] = |(datain[119:116] ^ 2);
  assign w780[49] = |(datain[115:112] ^ 0);
  assign w780[50] = |(datain[111:108] ^ 2);
  assign w780[51] = |(datain[107:104] ^ 5);
  assign w780[52] = |(datain[103:100] ^ 2);
  assign w780[53] = |(datain[99:96] ^ 5);
  assign w780[54] = |(datain[95:92] ^ 6);
  assign w780[55] = |(datain[91:88] ^ 2);
  assign w780[56] = |(datain[87:84] ^ 2);
  assign w780[57] = |(datain[83:80] ^ 11);
  assign w780[58] = |(datain[79:76] ^ 2);
  assign w780[59] = |(datain[75:72] ^ 5);
  assign w780[60] = |(datain[71:68] ^ 3);
  assign w780[61] = |(datain[67:64] ^ 0);
  assign comp[780] = ~(|w780);
  wire [64-1:0] w781;
  assign w781[0] = |(datain[311:308] ^ 6);
  assign w781[1] = |(datain[307:304] ^ 15);
  assign w781[2] = |(datain[303:300] ^ 7);
  assign w781[3] = |(datain[299:296] ^ 2);
  assign w781[4] = |(datain[295:292] ^ 2);
  assign w781[5] = |(datain[291:288] ^ 0);
  assign w781[6] = |(datain[287:284] ^ 2);
  assign w781[7] = |(datain[283:280] ^ 5);
  assign w781[8] = |(datain[279:276] ^ 2);
  assign w781[9] = |(datain[275:272] ^ 5);
  assign w781[10] = |(datain[271:268] ^ 6);
  assign w781[11] = |(datain[267:264] ^ 2);
  assign w781[12] = |(datain[263:260] ^ 2);
  assign w781[13] = |(datain[259:256] ^ 0);
  assign w781[14] = |(datain[255:252] ^ 6);
  assign w781[15] = |(datain[251:248] ^ 9);
  assign w781[16] = |(datain[247:244] ^ 6);
  assign w781[17] = |(datain[243:240] ^ 14);
  assign w781[18] = |(datain[239:236] ^ 2);
  assign w781[19] = |(datain[235:232] ^ 0);
  assign w781[20] = |(datain[231:228] ^ 2);
  assign w781[21] = |(datain[227:224] ^ 8);
  assign w781[22] = |(datain[223:220] ^ 2);
  assign w781[23] = |(datain[219:216] ^ 10);
  assign w781[24] = |(datain[215:212] ^ 2);
  assign w781[25] = |(datain[211:208] ^ 14);
  assign w781[26] = |(datain[207:204] ^ 6);
  assign w781[27] = |(datain[203:200] ^ 2);
  assign w781[28] = |(datain[199:196] ^ 6);
  assign w781[29] = |(datain[195:192] ^ 1);
  assign w781[30] = |(datain[191:188] ^ 7);
  assign w781[31] = |(datain[187:184] ^ 4);
  assign w781[32] = |(datain[183:180] ^ 2);
  assign w781[33] = |(datain[179:176] ^ 9);
  assign w781[34] = |(datain[175:172] ^ 2);
  assign w781[35] = |(datain[171:168] ^ 0);
  assign w781[36] = |(datain[167:164] ^ 6);
  assign w781[37] = |(datain[163:160] ^ 4);
  assign w781[38] = |(datain[159:156] ^ 6);
  assign w781[39] = |(datain[155:152] ^ 15);
  assign w781[40] = |(datain[151:148] ^ 2);
  assign w781[41] = |(datain[147:144] ^ 0);
  assign w781[42] = |(datain[143:140] ^ 6);
  assign w781[43] = |(datain[139:136] ^ 3);
  assign w781[44] = |(datain[135:132] ^ 6);
  assign w781[45] = |(datain[131:128] ^ 15);
  assign w781[46] = |(datain[127:124] ^ 7);
  assign w781[47] = |(datain[123:120] ^ 0);
  assign w781[48] = |(datain[119:116] ^ 7);
  assign w781[49] = |(datain[115:112] ^ 9);
  assign w781[50] = |(datain[111:108] ^ 2);
  assign w781[51] = |(datain[107:104] ^ 0);
  assign w781[52] = |(datain[103:100] ^ 2);
  assign w781[53] = |(datain[99:96] ^ 5);
  assign w781[54] = |(datain[95:92] ^ 3);
  assign w781[55] = |(datain[91:88] ^ 0);
  assign w781[56] = |(datain[87:84] ^ 2);
  assign w781[57] = |(datain[83:80] ^ 0);
  assign w781[58] = |(datain[79:76] ^ 2);
  assign w781[59] = |(datain[75:72] ^ 5);
  assign w781[60] = |(datain[71:68] ^ 2);
  assign w781[61] = |(datain[67:64] ^ 5);
  assign w781[62] = |(datain[63:60] ^ 6);
  assign w781[63] = |(datain[59:56] ^ 2);
  assign comp[781] = ~(|w781);
  wire [60-1:0] w782;
  assign w782[0] = |(datain[311:308] ^ 6);
  assign w782[1] = |(datain[307:304] ^ 15);
  assign w782[2] = |(datain[303:300] ^ 7);
  assign w782[3] = |(datain[299:296] ^ 2);
  assign w782[4] = |(datain[295:292] ^ 2);
  assign w782[5] = |(datain[291:288] ^ 0);
  assign w782[6] = |(datain[287:284] ^ 2);
  assign w782[7] = |(datain[283:280] ^ 5);
  assign w782[8] = |(datain[279:276] ^ 2);
  assign w782[9] = |(datain[275:272] ^ 5);
  assign w782[10] = |(datain[271:268] ^ 6);
  assign w782[11] = |(datain[267:264] ^ 2);
  assign w782[12] = |(datain[263:260] ^ 2);
  assign w782[13] = |(datain[259:256] ^ 0);
  assign w782[14] = |(datain[255:252] ^ 6);
  assign w782[15] = |(datain[251:248] ^ 9);
  assign w782[16] = |(datain[247:244] ^ 6);
  assign w782[17] = |(datain[243:240] ^ 14);
  assign w782[18] = |(datain[239:236] ^ 2);
  assign w782[19] = |(datain[235:232] ^ 0);
  assign w782[20] = |(datain[231:228] ^ 2);
  assign w782[21] = |(datain[227:224] ^ 8);
  assign w782[22] = |(datain[223:220] ^ 2);
  assign w782[23] = |(datain[219:216] ^ 10);
  assign w782[24] = |(datain[215:212] ^ 2);
  assign w782[25] = |(datain[211:208] ^ 14);
  assign w782[26] = |(datain[207:204] ^ 2);
  assign w782[27] = |(datain[203:200] ^ 10);
  assign w782[28] = |(datain[199:196] ^ 2);
  assign w782[29] = |(datain[195:192] ^ 9);
  assign w782[30] = |(datain[191:188] ^ 2);
  assign w782[31] = |(datain[187:184] ^ 0);
  assign w782[32] = |(datain[183:180] ^ 6);
  assign w782[33] = |(datain[179:176] ^ 4);
  assign w782[34] = |(datain[175:172] ^ 6);
  assign w782[35] = |(datain[171:168] ^ 15);
  assign w782[36] = |(datain[167:164] ^ 2);
  assign w782[37] = |(datain[163:160] ^ 0);
  assign w782[38] = |(datain[159:156] ^ 6);
  assign w782[39] = |(datain[155:152] ^ 3);
  assign w782[40] = |(datain[151:148] ^ 6);
  assign w782[41] = |(datain[147:144] ^ 15);
  assign w782[42] = |(datain[143:140] ^ 7);
  assign w782[43] = |(datain[139:136] ^ 0);
  assign w782[44] = |(datain[135:132] ^ 7);
  assign w782[45] = |(datain[131:128] ^ 9);
  assign w782[46] = |(datain[127:124] ^ 2);
  assign w782[47] = |(datain[123:120] ^ 0);
  assign w782[48] = |(datain[119:116] ^ 2);
  assign w782[49] = |(datain[115:112] ^ 5);
  assign w782[50] = |(datain[111:108] ^ 3);
  assign w782[51] = |(datain[107:104] ^ 0);
  assign w782[52] = |(datain[103:100] ^ 2);
  assign w782[53] = |(datain[99:96] ^ 0);
  assign w782[54] = |(datain[95:92] ^ 2);
  assign w782[55] = |(datain[91:88] ^ 5);
  assign w782[56] = |(datain[87:84] ^ 2);
  assign w782[57] = |(datain[83:80] ^ 5);
  assign w782[58] = |(datain[79:76] ^ 6);
  assign w782[59] = |(datain[75:72] ^ 2);
  assign comp[782] = ~(|w782);
  wire [66-1:0] w783;
  assign w783[0] = |(datain[311:308] ^ 6);
  assign w783[1] = |(datain[307:304] ^ 6);
  assign w783[2] = |(datain[303:300] ^ 6);
  assign w783[3] = |(datain[299:296] ^ 15);
  assign w783[4] = |(datain[295:292] ^ 7);
  assign w783[5] = |(datain[291:288] ^ 2);
  assign w783[6] = |(datain[287:284] ^ 2);
  assign w783[7] = |(datain[283:280] ^ 0);
  assign w783[8] = |(datain[279:276] ^ 2);
  assign w783[9] = |(datain[275:272] ^ 5);
  assign w783[10] = |(datain[271:268] ^ 2);
  assign w783[11] = |(datain[267:264] ^ 5);
  assign w783[12] = |(datain[263:260] ^ 6);
  assign w783[13] = |(datain[259:256] ^ 2);
  assign w783[14] = |(datain[255:252] ^ 2);
  assign w783[15] = |(datain[251:248] ^ 0);
  assign w783[16] = |(datain[247:244] ^ 6);
  assign w783[17] = |(datain[243:240] ^ 9);
  assign w783[18] = |(datain[239:236] ^ 6);
  assign w783[19] = |(datain[235:232] ^ 14);
  assign w783[20] = |(datain[231:228] ^ 2);
  assign w783[21] = |(datain[227:224] ^ 0);
  assign w783[22] = |(datain[223:220] ^ 2);
  assign w783[23] = |(datain[219:216] ^ 8);
  assign w783[24] = |(datain[215:212] ^ 2);
  assign w783[25] = |(datain[211:208] ^ 10);
  assign w783[26] = |(datain[207:204] ^ 2);
  assign w783[27] = |(datain[203:200] ^ 14);
  assign w783[28] = |(datain[199:196] ^ 6);
  assign w783[29] = |(datain[195:192] ^ 2);
  assign w783[30] = |(datain[191:188] ^ 6);
  assign w783[31] = |(datain[187:184] ^ 1);
  assign w783[32] = |(datain[183:180] ^ 7);
  assign w783[33] = |(datain[179:176] ^ 4);
  assign w783[34] = |(datain[175:172] ^ 2);
  assign w783[35] = |(datain[171:168] ^ 9);
  assign w783[36] = |(datain[167:164] ^ 2);
  assign w783[37] = |(datain[163:160] ^ 0);
  assign w783[38] = |(datain[159:156] ^ 6);
  assign w783[39] = |(datain[155:152] ^ 4);
  assign w783[40] = |(datain[151:148] ^ 6);
  assign w783[41] = |(datain[147:144] ^ 15);
  assign w783[42] = |(datain[143:140] ^ 2);
  assign w783[43] = |(datain[139:136] ^ 0);
  assign w783[44] = |(datain[135:132] ^ 6);
  assign w783[45] = |(datain[131:128] ^ 3);
  assign w783[46] = |(datain[127:124] ^ 6);
  assign w783[47] = |(datain[123:120] ^ 15);
  assign w783[48] = |(datain[119:116] ^ 7);
  assign w783[49] = |(datain[115:112] ^ 0);
  assign w783[50] = |(datain[111:108] ^ 7);
  assign w783[51] = |(datain[107:104] ^ 9);
  assign w783[52] = |(datain[103:100] ^ 2);
  assign w783[53] = |(datain[99:96] ^ 0);
  assign w783[54] = |(datain[95:92] ^ 2);
  assign w783[55] = |(datain[91:88] ^ 5);
  assign w783[56] = |(datain[87:84] ^ 3);
  assign w783[57] = |(datain[83:80] ^ 0);
  assign w783[58] = |(datain[79:76] ^ 2);
  assign w783[59] = |(datain[75:72] ^ 0);
  assign w783[60] = |(datain[71:68] ^ 2);
  assign w783[61] = |(datain[67:64] ^ 5);
  assign w783[62] = |(datain[63:60] ^ 6);
  assign w783[63] = |(datain[59:56] ^ 1);
  assign w783[64] = |(datain[55:52] ^ 2);
  assign w783[65] = |(datain[51:48] ^ 5);
  assign comp[783] = ~(|w783);
  wire [60-1:0] w784;
  assign w784[0] = |(datain[311:308] ^ 6);
  assign w784[1] = |(datain[307:304] ^ 15);
  assign w784[2] = |(datain[303:300] ^ 7);
  assign w784[3] = |(datain[299:296] ^ 2);
  assign w784[4] = |(datain[295:292] ^ 2);
  assign w784[5] = |(datain[291:288] ^ 0);
  assign w784[6] = |(datain[287:284] ^ 2);
  assign w784[7] = |(datain[283:280] ^ 5);
  assign w784[8] = |(datain[279:276] ^ 2);
  assign w784[9] = |(datain[275:272] ^ 5);
  assign w784[10] = |(datain[271:268] ^ 6);
  assign w784[11] = |(datain[267:264] ^ 2);
  assign w784[12] = |(datain[263:260] ^ 2);
  assign w784[13] = |(datain[259:256] ^ 0);
  assign w784[14] = |(datain[255:252] ^ 6);
  assign w784[15] = |(datain[251:248] ^ 9);
  assign w784[16] = |(datain[247:244] ^ 6);
  assign w784[17] = |(datain[243:240] ^ 14);
  assign w784[18] = |(datain[239:236] ^ 2);
  assign w784[19] = |(datain[235:232] ^ 0);
  assign w784[20] = |(datain[231:228] ^ 2);
  assign w784[21] = |(datain[227:224] ^ 8);
  assign w784[22] = |(datain[223:220] ^ 2);
  assign w784[23] = |(datain[219:216] ^ 10);
  assign w784[24] = |(datain[215:212] ^ 2);
  assign w784[25] = |(datain[211:208] ^ 14);
  assign w784[26] = |(datain[207:204] ^ 2);
  assign w784[27] = |(datain[203:200] ^ 10);
  assign w784[28] = |(datain[199:196] ^ 2);
  assign w784[29] = |(datain[195:192] ^ 9);
  assign w784[30] = |(datain[191:188] ^ 2);
  assign w784[31] = |(datain[187:184] ^ 0);
  assign w784[32] = |(datain[183:180] ^ 6);
  assign w784[33] = |(datain[179:176] ^ 4);
  assign w784[34] = |(datain[175:172] ^ 6);
  assign w784[35] = |(datain[171:168] ^ 15);
  assign w784[36] = |(datain[167:164] ^ 2);
  assign w784[37] = |(datain[163:160] ^ 0);
  assign w784[38] = |(datain[159:156] ^ 6);
  assign w784[39] = |(datain[155:152] ^ 3);
  assign w784[40] = |(datain[151:148] ^ 6);
  assign w784[41] = |(datain[147:144] ^ 15);
  assign w784[42] = |(datain[143:140] ^ 7);
  assign w784[43] = |(datain[139:136] ^ 0);
  assign w784[44] = |(datain[135:132] ^ 7);
  assign w784[45] = |(datain[131:128] ^ 9);
  assign w784[46] = |(datain[127:124] ^ 2);
  assign w784[47] = |(datain[123:120] ^ 0);
  assign w784[48] = |(datain[119:116] ^ 2);
  assign w784[49] = |(datain[115:112] ^ 5);
  assign w784[50] = |(datain[111:108] ^ 2);
  assign w784[51] = |(datain[107:104] ^ 5);
  assign w784[52] = |(datain[103:100] ^ 6);
  assign w784[53] = |(datain[99:96] ^ 2);
  assign w784[54] = |(datain[95:92] ^ 2);
  assign w784[55] = |(datain[91:88] ^ 11);
  assign w784[56] = |(datain[87:84] ^ 2);
  assign w784[57] = |(datain[83:80] ^ 5);
  assign w784[58] = |(datain[79:76] ^ 3);
  assign w784[59] = |(datain[75:72] ^ 0);
  assign comp[784] = ~(|w784);
  wire [52-1:0] w785;
  assign w785[0] = |(datain[311:308] ^ 7);
  assign w785[1] = |(datain[307:304] ^ 10);
  assign w785[2] = |(datain[303:300] ^ 3);
  assign w785[3] = |(datain[299:296] ^ 11);
  assign w785[4] = |(datain[295:292] ^ 12);
  assign w785[5] = |(datain[291:288] ^ 14);
  assign w785[6] = |(datain[287:284] ^ 0);
  assign w785[7] = |(datain[283:280] ^ 4);
  assign w785[8] = |(datain[279:276] ^ 11);
  assign w785[9] = |(datain[275:272] ^ 11);
  assign w785[10] = |(datain[271:268] ^ 0);
  assign w785[11] = |(datain[267:264] ^ 3);
  assign w785[12] = |(datain[263:260] ^ 0);
  assign w785[13] = |(datain[259:256] ^ 1);
  assign w785[14] = |(datain[255:252] ^ 11);
  assign w785[15] = |(datain[251:248] ^ 8);
  assign w785[16] = |(datain[247:244] ^ 10);
  assign w785[17] = |(datain[243:240] ^ 6);
  assign w785[18] = |(datain[239:236] ^ 0);
  assign w785[19] = |(datain[235:232] ^ 4);
  assign w785[20] = |(datain[231:228] ^ 8);
  assign w785[21] = |(datain[227:224] ^ 11);
  assign w785[22] = |(datain[223:220] ^ 0);
  assign w785[23] = |(datain[219:216] ^ 14);
  assign w785[24] = |(datain[215:212] ^ 10);
  assign w785[25] = |(datain[211:208] ^ 11);
  assign w785[26] = |(datain[207:204] ^ 0);
  assign w785[27] = |(datain[203:200] ^ 4);
  assign w785[28] = |(datain[199:196] ^ 3);
  assign w785[29] = |(datain[195:192] ^ 1);
  assign w785[30] = |(datain[191:188] ^ 0);
  assign w785[31] = |(datain[187:184] ^ 15);
  assign w785[32] = |(datain[183:180] ^ 4);
  assign w785[33] = |(datain[179:176] ^ 3);
  assign w785[34] = |(datain[175:172] ^ 4);
  assign w785[35] = |(datain[171:168] ^ 3);
  assign w785[36] = |(datain[167:164] ^ 3);
  assign w785[37] = |(datain[163:160] ^ 11);
  assign w785[38] = |(datain[159:156] ^ 13);
  assign w785[39] = |(datain[155:152] ^ 8);
  assign w785[40] = |(datain[151:148] ^ 7);
  assign w785[41] = |(datain[147:144] ^ 6);
  assign w785[42] = |(datain[143:140] ^ 15);
  assign w785[43] = |(datain[139:136] ^ 8);
  assign w785[44] = |(datain[135:132] ^ 12);
  assign w785[45] = |(datain[131:128] ^ 3);
  assign w785[46] = |(datain[127:124] ^ 14);
  assign w785[47] = |(datain[123:120] ^ 8);
  assign w785[48] = |(datain[119:116] ^ 14);
  assign w785[49] = |(datain[115:112] ^ 10);
  assign w785[50] = |(datain[111:108] ^ 15);
  assign w785[51] = |(datain[107:104] ^ 15);
  assign comp[785] = ~(|w785);
  wire [44-1:0] w786;
  assign w786[0] = |(datain[311:308] ^ 0);
  assign w786[1] = |(datain[307:304] ^ 1);
  assign w786[2] = |(datain[303:300] ^ 0);
  assign w786[3] = |(datain[299:296] ^ 1);
  assign w786[4] = |(datain[295:292] ^ 8);
  assign w786[5] = |(datain[291:288] ^ 1);
  assign w786[6] = |(datain[287:284] ^ 12);
  assign w786[7] = |(datain[283:280] ^ 7);
  assign w786[8] = |(datain[279:276] ^ 0);
  assign w786[9] = |(datain[275:272] ^ 0);
  assign w786[10] = |(datain[271:268] ^ 0);
  assign w786[11] = |(datain[267:264] ^ 1);
  assign w786[12] = |(datain[263:260] ^ 14);
  assign w786[13] = |(datain[259:256] ^ 8);
  assign w786[14] = |(datain[255:252] ^ 0);
  assign w786[15] = |(datain[251:248] ^ 3);
  assign w786[16] = |(datain[247:244] ^ 0);
  assign w786[17] = |(datain[243:240] ^ 0);
  assign w786[18] = |(datain[239:236] ^ 14);
  assign w786[19] = |(datain[235:232] ^ 9);
  assign w786[20] = |(datain[231:228] ^ 3);
  assign w786[21] = |(datain[227:224] ^ 9);
  assign w786[22] = |(datain[223:220] ^ 0);
  assign w786[23] = |(datain[219:216] ^ 2);
  assign w786[24] = |(datain[215:212] ^ 11);
  assign w786[25] = |(datain[211:208] ^ 9);
  assign w786[26] = |(datain[207:204] ^ 3);
  assign w786[27] = |(datain[203:200] ^ 14);
  assign w786[28] = |(datain[199:196] ^ 0);
  assign w786[29] = |(datain[195:192] ^ 5);
  assign w786[30] = |(datain[191:188] ^ 11);
  assign w786[31] = |(datain[187:184] ^ 11);
  assign w786[32] = |(datain[183:180] ^ 5);
  assign w786[33] = |(datain[179:176] ^ 3);
  assign w786[34] = |(datain[175:172] ^ 0);
  assign w786[35] = |(datain[171:168] ^ 2);
  assign w786[36] = |(datain[167:164] ^ 0);
  assign w786[37] = |(datain[163:160] ^ 3);
  assign w786[38] = |(datain[159:156] ^ 13);
  assign w786[39] = |(datain[155:152] ^ 15);
  assign w786[40] = |(datain[151:148] ^ 8);
  assign w786[41] = |(datain[147:144] ^ 0);
  assign w786[42] = |(datain[143:140] ^ 3);
  assign w786[43] = |(datain[139:136] ^ 7);
  assign comp[786] = ~(|w786);
  wire [30-1:0] w787;
  assign w787[0] = |(datain[311:308] ^ 7);
  assign w787[1] = |(datain[307:304] ^ 3);
  assign w787[2] = |(datain[303:300] ^ 0);
  assign w787[3] = |(datain[299:296] ^ 3);
  assign w787[4] = |(datain[295:292] ^ 11);
  assign w787[5] = |(datain[291:288] ^ 14);
  assign w787[6] = |(datain[287:284] ^ 3);
  assign w787[7] = |(datain[283:280] ^ 9);
  assign w787[8] = |(datain[279:276] ^ 0);
  assign w787[9] = |(datain[275:272] ^ 1);
  assign w787[10] = |(datain[271:268] ^ 8);
  assign w787[11] = |(datain[267:264] ^ 11);
  assign w787[12] = |(datain[263:260] ^ 15);
  assign w787[13] = |(datain[259:256] ^ 14);
  assign w787[14] = |(datain[255:252] ^ 15);
  assign w787[15] = |(datain[251:248] ^ 12);
  assign w787[16] = |(datain[247:244] ^ 10);
  assign w787[17] = |(datain[243:240] ^ 13);
  assign w787[18] = |(datain[239:236] ^ 3);
  assign w787[19] = |(datain[235:232] ^ 3);
  assign w787[20] = |(datain[231:228] ^ 0);
  assign w787[21] = |(datain[227:224] ^ 6);
  assign w787[22] = |(datain[223:220] ^ 0);
  assign w787[23] = |(datain[219:216] ^ 3);
  assign w787[24] = |(datain[215:212] ^ 0);
  assign w787[25] = |(datain[211:208] ^ 1);
  assign w787[26] = |(datain[207:204] ^ 10);
  assign w787[27] = |(datain[203:200] ^ 11);
  assign w787[28] = |(datain[199:196] ^ 4);
  assign w787[29] = |(datain[195:192] ^ 9);
  assign comp[787] = ~(|w787);
  wire [42-1:0] w788;
  assign w788[0] = |(datain[311:308] ^ 0);
  assign w788[1] = |(datain[307:304] ^ 15);
  assign w788[2] = |(datain[303:300] ^ 0);
  assign w788[3] = |(datain[299:296] ^ 1);
  assign w788[4] = |(datain[295:292] ^ 8);
  assign w788[5] = |(datain[291:288] ^ 10);
  assign w788[6] = |(datain[287:284] ^ 2);
  assign w788[7] = |(datain[283:280] ^ 6);
  assign w788[8] = |(datain[279:276] ^ 0);
  assign w788[9] = |(datain[275:272] ^ 14);
  assign w788[10] = |(datain[271:268] ^ 0);
  assign w788[11] = |(datain[267:264] ^ 1);
  assign w788[12] = |(datain[263:260] ^ 11);
  assign w788[13] = |(datain[259:256] ^ 9);
  assign w788[14] = |(datain[255:252] ^ 5);
  assign w788[15] = |(datain[251:248] ^ 3);
  assign w788[16] = |(datain[247:244] ^ 0);
  assign w788[17] = |(datain[243:240] ^ 2);
  assign w788[18] = |(datain[239:236] ^ 8);
  assign w788[19] = |(datain[235:232] ^ 10);
  assign w788[20] = |(datain[231:228] ^ 0);
  assign w788[21] = |(datain[227:224] ^ 4);
  assign w788[22] = |(datain[223:220] ^ 3);
  assign w788[23] = |(datain[219:216] ^ 2);
  assign w788[24] = |(datain[215:212] ^ 12);
  assign w788[25] = |(datain[211:208] ^ 4);
  assign w788[26] = |(datain[207:204] ^ 8);
  assign w788[27] = |(datain[203:200] ^ 8);
  assign w788[28] = |(datain[199:196] ^ 0);
  assign w788[29] = |(datain[195:192] ^ 4);
  assign w788[30] = |(datain[191:188] ^ 4);
  assign w788[31] = |(datain[187:184] ^ 6);
  assign w788[32] = |(datain[183:180] ^ 3);
  assign w788[33] = |(datain[179:176] ^ 11);
  assign w788[34] = |(datain[175:172] ^ 15);
  assign w788[35] = |(datain[171:168] ^ 1);
  assign w788[36] = |(datain[167:164] ^ 7);
  assign w788[37] = |(datain[163:160] ^ 5);
  assign w788[38] = |(datain[159:156] ^ 15);
  assign w788[39] = |(datain[155:152] ^ 5);
  assign w788[40] = |(datain[151:148] ^ 12);
  assign w788[41] = |(datain[147:144] ^ 3);
  assign comp[788] = ~(|w788);
  wire [44-1:0] w789;
  assign w789[0] = |(datain[311:308] ^ 12);
  assign w789[1] = |(datain[307:304] ^ 13);
  assign w789[2] = |(datain[303:300] ^ 2);
  assign w789[3] = |(datain[299:296] ^ 1);
  assign w789[4] = |(datain[295:292] ^ 11);
  assign w789[5] = |(datain[291:288] ^ 8);
  assign w789[6] = |(datain[287:284] ^ 2);
  assign w789[7] = |(datain[283:280] ^ 4);
  assign w789[8] = |(datain[279:276] ^ 2);
  assign w789[9] = |(datain[275:272] ^ 5);
  assign w789[10] = |(datain[271:268] ^ 5);
  assign w789[11] = |(datain[267:264] ^ 10);
  assign w789[12] = |(datain[263:260] ^ 1);
  assign w789[13] = |(datain[259:256] ^ 15);
  assign w789[14] = |(datain[255:252] ^ 12);
  assign w789[15] = |(datain[251:248] ^ 13);
  assign w789[16] = |(datain[247:244] ^ 2);
  assign w789[17] = |(datain[243:240] ^ 1);
  assign w789[18] = |(datain[239:236] ^ 0);
  assign w789[19] = |(datain[235:232] ^ 6);
  assign w789[20] = |(datain[231:228] ^ 1);
  assign w789[21] = |(datain[227:224] ^ 15);
  assign w789[22] = |(datain[223:220] ^ 11);
  assign w789[23] = |(datain[219:216] ^ 15);
  assign w789[24] = |(datain[215:212] ^ 0);
  assign w789[25] = |(datain[211:208] ^ 0);
  assign w789[26] = |(datain[207:204] ^ 0);
  assign w789[27] = |(datain[203:200] ^ 1);
  assign w789[28] = |(datain[199:196] ^ 5);
  assign w789[29] = |(datain[195:192] ^ 7);
  assign w789[30] = |(datain[191:188] ^ 12);
  assign w789[31] = |(datain[187:184] ^ 2);
  assign w789[32] = |(datain[183:180] ^ 15);
  assign w789[33] = |(datain[179:176] ^ 15);
  assign w789[34] = |(datain[175:172] ^ 15);
  assign w789[35] = |(datain[171:168] ^ 15);
  assign w789[36] = |(datain[167:164] ^ 11);
  assign w789[37] = |(datain[163:160] ^ 4);
  assign w789[38] = |(datain[159:156] ^ 4);
  assign w789[39] = |(datain[155:152] ^ 15);
  assign w789[40] = |(datain[151:148] ^ 12);
  assign w789[41] = |(datain[147:144] ^ 13);
  assign w789[42] = |(datain[143:140] ^ 2);
  assign w789[43] = |(datain[139:136] ^ 1);
  assign comp[789] = ~(|w789);
  wire [28-1:0] w790;
  assign w790[0] = |(datain[311:308] ^ 7);
  assign w790[1] = |(datain[307:304] ^ 4);
  assign w790[2] = |(datain[303:300] ^ 2);
  assign w790[3] = |(datain[299:296] ^ 0);
  assign w790[4] = |(datain[295:292] ^ 5);
  assign w790[5] = |(datain[291:288] ^ 0);
  assign w790[6] = |(datain[287:284] ^ 3);
  assign w790[7] = |(datain[283:280] ^ 13);
  assign w790[8] = |(datain[279:276] ^ 0);
  assign w790[9] = |(datain[275:272] ^ 0);
  assign w790[10] = |(datain[271:268] ^ 5);
  assign w790[11] = |(datain[267:264] ^ 7);
  assign w790[12] = |(datain[263:260] ^ 7);
  assign w790[13] = |(datain[259:256] ^ 4);
  assign w790[14] = |(datain[255:252] ^ 13);
  assign w790[15] = |(datain[251:248] ^ 7);
  assign w790[16] = |(datain[247:244] ^ 8);
  assign w790[17] = |(datain[243:240] ^ 0);
  assign w790[18] = |(datain[239:236] ^ 15);
  assign w790[19] = |(datain[235:232] ^ 12);
  assign w790[20] = |(datain[231:228] ^ 3);
  assign w790[21] = |(datain[227:224] ^ 15);
  assign w790[22] = |(datain[223:220] ^ 7);
  assign w790[23] = |(datain[219:216] ^ 4);
  assign w790[24] = |(datain[215:212] ^ 9);
  assign w790[25] = |(datain[211:208] ^ 10);
  assign w790[26] = |(datain[207:204] ^ 5);
  assign w790[27] = |(datain[203:200] ^ 3);
  assign comp[790] = ~(|w790);
  wire [32-1:0] w791;
  assign w791[0] = |(datain[311:308] ^ 0);
  assign w791[1] = |(datain[307:304] ^ 1);
  assign w791[2] = |(datain[303:300] ^ 3);
  assign w791[3] = |(datain[299:296] ^ 11);
  assign w791[4] = |(datain[295:292] ^ 3);
  assign w791[5] = |(datain[291:288] ^ 6);
  assign w791[6] = |(datain[287:284] ^ 15);
  assign w791[7] = |(datain[283:280] ^ 14);
  assign w791[8] = |(datain[279:276] ^ 0);
  assign w791[9] = |(datain[275:272] ^ 2);
  assign w791[10] = |(datain[271:268] ^ 7);
  assign w791[11] = |(datain[267:264] ^ 5);
  assign w791[12] = |(datain[263:260] ^ 0);
  assign w791[13] = |(datain[259:256] ^ 2);
  assign w791[14] = |(datain[255:252] ^ 11);
  assign w791[15] = |(datain[251:248] ^ 4);
  assign w791[16] = |(datain[247:244] ^ 3);
  assign w791[17] = |(datain[243:240] ^ 15);
  assign w791[18] = |(datain[239:236] ^ 14);
  assign w791[19] = |(datain[235:232] ^ 9);
  assign w791[20] = |(datain[231:228] ^ 10);
  assign w791[21] = |(datain[227:224] ^ 1);
  assign w791[22] = |(datain[223:220] ^ 15);
  assign w791[23] = |(datain[219:216] ^ 14);
  assign w791[24] = |(datain[215:212] ^ 5);
  assign w791[25] = |(datain[211:208] ^ 3);
  assign w791[26] = |(datain[207:204] ^ 11);
  assign w791[27] = |(datain[203:200] ^ 8);
  assign w791[28] = |(datain[199:196] ^ 2);
  assign w791[29] = |(datain[195:192] ^ 0);
  assign w791[30] = |(datain[191:188] ^ 1);
  assign w791[31] = |(datain[187:184] ^ 2);
  assign comp[791] = ~(|w791);
  wire [32-1:0] w792;
  assign w792[0] = |(datain[311:308] ^ 12);
  assign w792[1] = |(datain[307:304] ^ 13);
  assign w792[2] = |(datain[303:300] ^ 2);
  assign w792[3] = |(datain[299:296] ^ 1);
  assign w792[4] = |(datain[295:292] ^ 7);
  assign w792[5] = |(datain[291:288] ^ 2);
  assign w792[6] = |(datain[287:284] ^ 0);
  assign w792[7] = |(datain[283:280] ^ 12);
  assign w792[8] = |(datain[279:276] ^ 11);
  assign w792[9] = |(datain[275:272] ^ 4);
  assign w792[10] = |(datain[271:268] ^ 4);
  assign w792[11] = |(datain[267:264] ^ 0);
  assign w792[12] = |(datain[263:260] ^ 11);
  assign w792[13] = |(datain[259:256] ^ 9);
  assign w792[14] = |(datain[255:252] ^ 0);
  assign w792[15] = |(datain[251:248] ^ 3);
  assign w792[16] = |(datain[247:244] ^ 0);
  assign w792[17] = |(datain[243:240] ^ 0);
  assign w792[18] = |(datain[239:236] ^ 11);
  assign w792[19] = |(datain[235:232] ^ 10);
  assign w792[20] = |(datain[231:228] ^ 4);
  assign w792[21] = |(datain[227:224] ^ 7);
  assign w792[22] = |(datain[223:220] ^ 0);
  assign w792[23] = |(datain[219:216] ^ 0);
  assign w792[24] = |(datain[215:212] ^ 0);
  assign w792[25] = |(datain[211:208] ^ 3);
  assign w792[26] = |(datain[207:204] ^ 13);
  assign w792[27] = |(datain[203:200] ^ 6);
  assign w792[28] = |(datain[199:196] ^ 12);
  assign w792[29] = |(datain[195:192] ^ 13);
  assign w792[30] = |(datain[191:188] ^ 2);
  assign w792[31] = |(datain[187:184] ^ 1);
  assign comp[792] = ~(|w792);
  wire [50-1:0] w793;
  assign w793[0] = |(datain[311:308] ^ 4);
  assign w793[1] = |(datain[307:304] ^ 4);
  assign w793[2] = |(datain[303:300] ^ 11);
  assign w793[3] = |(datain[299:296] ^ 11);
  assign w793[4] = |(datain[295:292] ^ 5);
  assign w793[5] = |(datain[291:288] ^ 12);
  assign w793[6] = |(datain[287:284] ^ 7);
  assign w793[7] = |(datain[283:280] ^ 12);
  assign w793[8] = |(datain[279:276] ^ 11);
  assign w793[9] = |(datain[275:272] ^ 14);
  assign w793[10] = |(datain[271:268] ^ 0);
  assign w793[11] = |(datain[267:264] ^ 4);
  assign w793[12] = |(datain[263:260] ^ 0);
  assign w793[13] = |(datain[259:256] ^ 1);
  assign w793[14] = |(datain[255:252] ^ 8);
  assign w793[15] = |(datain[251:248] ^ 10);
  assign w793[16] = |(datain[247:244] ^ 0);
  assign w793[17] = |(datain[243:240] ^ 7);
  assign w793[18] = |(datain[239:236] ^ 3);
  assign w793[19] = |(datain[235:232] ^ 4);
  assign w793[20] = |(datain[231:228] ^ 9);
  assign w793[21] = |(datain[227:224] ^ 0);
  assign w793[22] = |(datain[223:220] ^ 4);
  assign w793[23] = |(datain[219:216] ^ 14);
  assign w793[24] = |(datain[215:212] ^ 3);
  assign w793[25] = |(datain[211:208] ^ 0);
  assign w793[26] = |(datain[207:204] ^ 0);
  assign w793[27] = |(datain[203:200] ^ 0);
  assign w793[28] = |(datain[199:196] ^ 0);
  assign w793[29] = |(datain[195:192] ^ 11);
  assign w793[30] = |(datain[191:188] ^ 15);
  assign w793[31] = |(datain[187:184] ^ 6);
  assign w793[32] = |(datain[183:180] ^ 7);
  assign w793[33] = |(datain[179:176] ^ 5);
  assign w793[34] = |(datain[175:172] ^ 15);
  assign w793[35] = |(datain[171:168] ^ 9);
  assign w793[36] = |(datain[167:164] ^ 12);
  assign w793[37] = |(datain[163:160] ^ 3);
  assign w793[38] = |(datain[159:156] ^ 1);
  assign w793[39] = |(datain[155:152] ^ 4);
  assign w793[40] = |(datain[151:148] ^ 9);
  assign w793[41] = |(datain[147:144] ^ 10);
  assign w793[42] = |(datain[143:140] ^ 0);
  assign w793[43] = |(datain[139:136] ^ 0);
  assign w793[44] = |(datain[135:132] ^ 15);
  assign w793[45] = |(datain[131:128] ^ 0);
  assign w793[46] = |(datain[127:124] ^ 0);
  assign w793[47] = |(datain[123:120] ^ 0);
  assign w793[48] = |(datain[119:116] ^ 7);
  assign w793[49] = |(datain[115:112] ^ 12);
  assign comp[793] = ~(|w793);
  wire [44-1:0] w794;
  assign w794[0] = |(datain[311:308] ^ 7);
  assign w794[1] = |(datain[307:304] ^ 12);
  assign w794[2] = |(datain[303:300] ^ 11);
  assign w794[3] = |(datain[299:296] ^ 14);
  assign w794[4] = |(datain[295:292] ^ 15);
  assign w794[5] = |(datain[291:288] ^ 14);
  assign w794[6] = |(datain[287:284] ^ 0);
  assign w794[7] = |(datain[283:280] ^ 0);
  assign w794[8] = |(datain[279:276] ^ 8);
  assign w794[9] = |(datain[275:272] ^ 10);
  assign w794[10] = |(datain[271:268] ^ 0);
  assign w794[11] = |(datain[267:264] ^ 7);
  assign w794[12] = |(datain[263:260] ^ 3);
  assign w794[13] = |(datain[259:256] ^ 4);
  assign w794[14] = |(datain[255:252] ^ 9);
  assign w794[15] = |(datain[251:248] ^ 0);
  assign w794[16] = |(datain[247:244] ^ 4);
  assign w794[17] = |(datain[243:240] ^ 14);
  assign w794[18] = |(datain[239:236] ^ 3);
  assign w794[19] = |(datain[235:232] ^ 0);
  assign w794[20] = |(datain[231:228] ^ 0);
  assign w794[21] = |(datain[227:224] ^ 0);
  assign w794[22] = |(datain[223:220] ^ 0);
  assign w794[23] = |(datain[219:216] ^ 11);
  assign w794[24] = |(datain[215:212] ^ 15);
  assign w794[25] = |(datain[211:208] ^ 6);
  assign w794[26] = |(datain[207:204] ^ 7);
  assign w794[27] = |(datain[203:200] ^ 5);
  assign w794[28] = |(datain[199:196] ^ 15);
  assign w794[29] = |(datain[195:192] ^ 9);
  assign w794[30] = |(datain[191:188] ^ 12);
  assign w794[31] = |(datain[187:184] ^ 3);
  assign w794[32] = |(datain[183:180] ^ 4);
  assign w794[33] = |(datain[179:176] ^ 4);
  assign w794[34] = |(datain[175:172] ^ 10);
  assign w794[35] = |(datain[171:168] ^ 13);
  assign w794[36] = |(datain[167:164] ^ 0);
  assign w794[37] = |(datain[163:160] ^ 0);
  assign w794[38] = |(datain[159:156] ^ 15);
  assign w794[39] = |(datain[155:152] ^ 0);
  assign w794[40] = |(datain[151:148] ^ 0);
  assign w794[41] = |(datain[147:144] ^ 0);
  assign w794[42] = |(datain[143:140] ^ 7);
  assign w794[43] = |(datain[139:136] ^ 2);
  assign comp[794] = ~(|w794);
  wire [76-1:0] w795;
  assign w795[0] = |(datain[311:308] ^ 15);
  assign w795[1] = |(datain[307:304] ^ 14);
  assign w795[2] = |(datain[303:300] ^ 11);
  assign w795[3] = |(datain[299:296] ^ 9);
  assign w795[4] = |(datain[295:292] ^ 0);
  assign w795[5] = |(datain[291:288] ^ 0);
  assign w795[6] = |(datain[287:284] ^ 0);
  assign w795[7] = |(datain[283:280] ^ 2);
  assign w795[8] = |(datain[279:276] ^ 15);
  assign w795[9] = |(datain[275:272] ^ 7);
  assign w795[10] = |(datain[271:268] ^ 15);
  assign w795[11] = |(datain[267:264] ^ 1);
  assign w795[12] = |(datain[263:260] ^ 8);
  assign w795[13] = |(datain[259:256] ^ 3);
  assign w795[14] = |(datain[255:252] ^ 15);
  assign w795[15] = |(datain[251:248] ^ 10);
  assign w795[16] = |(datain[247:244] ^ 0);
  assign w795[17] = |(datain[243:240] ^ 0);
  assign w795[18] = |(datain[239:236] ^ 7);
  assign w795[19] = |(datain[235:232] ^ 4);
  assign w795[20] = |(datain[231:228] ^ 0);
  assign w795[21] = |(datain[227:224] ^ 1);
  assign w795[22] = |(datain[223:220] ^ 4);
  assign w795[23] = |(datain[219:216] ^ 0);
  assign w795[24] = |(datain[215:212] ^ 10);
  assign w795[25] = |(datain[211:208] ^ 3);
  assign w795[26] = |(datain[207:204] ^ 10);
  assign w795[27] = |(datain[203:200] ^ 3);
  assign w795[28] = |(datain[199:196] ^ 0);
  assign w795[29] = |(datain[195:192] ^ 2);
  assign w795[30] = |(datain[191:188] ^ 8);
  assign w795[31] = |(datain[187:184] ^ 9);
  assign w795[32] = |(datain[183:180] ^ 1);
  assign w795[33] = |(datain[179:176] ^ 6);
  assign w795[34] = |(datain[175:172] ^ 10);
  assign w795[35] = |(datain[171:168] ^ 1);
  assign w795[36] = |(datain[167:164] ^ 0);
  assign w795[37] = |(datain[163:160] ^ 2);
  assign w795[38] = |(datain[159:156] ^ 3);
  assign w795[39] = |(datain[155:152] ^ 3);
  assign w795[40] = |(datain[151:148] ^ 13);
  assign w795[41] = |(datain[147:144] ^ 2);
  assign w795[42] = |(datain[143:140] ^ 3);
  assign w795[43] = |(datain[139:136] ^ 3);
  assign w795[44] = |(datain[135:132] ^ 12);
  assign w795[45] = |(datain[131:128] ^ 9);
  assign w795[46] = |(datain[127:124] ^ 11);
  assign w795[47] = |(datain[123:120] ^ 8);
  assign w795[48] = |(datain[119:116] ^ 0);
  assign w795[49] = |(datain[115:112] ^ 0);
  assign w795[50] = |(datain[111:108] ^ 4);
  assign w795[51] = |(datain[107:104] ^ 2);
  assign w795[52] = |(datain[103:100] ^ 12);
  assign w795[53] = |(datain[99:96] ^ 13);
  assign w795[54] = |(datain[95:92] ^ 2);
  assign w795[55] = |(datain[91:88] ^ 1);
  assign w795[56] = |(datain[87:84] ^ 11);
  assign w795[57] = |(datain[83:80] ^ 9);
  assign w795[58] = |(datain[79:76] ^ 1);
  assign w795[59] = |(datain[75:72] ^ 12);
  assign w795[60] = |(datain[71:68] ^ 0);
  assign w795[61] = |(datain[67:64] ^ 0);
  assign w795[62] = |(datain[63:60] ^ 11);
  assign w795[63] = |(datain[59:56] ^ 10);
  assign w795[64] = |(datain[55:52] ^ 9);
  assign w795[65] = |(datain[51:48] ^ 15);
  assign w795[66] = |(datain[47:44] ^ 0);
  assign w795[67] = |(datain[43:40] ^ 2);
  assign w795[68] = |(datain[39:36] ^ 11);
  assign w795[69] = |(datain[35:32] ^ 4);
  assign w795[70] = |(datain[31:28] ^ 4);
  assign w795[71] = |(datain[27:24] ^ 0);
  assign w795[72] = |(datain[23:20] ^ 12);
  assign w795[73] = |(datain[19:16] ^ 13);
  assign w795[74] = |(datain[15:12] ^ 2);
  assign w795[75] = |(datain[11:8] ^ 1);
  assign comp[795] = ~(|w795);
  wire [32-1:0] w796;
  assign w796[0] = |(datain[311:308] ^ 1);
  assign w796[1] = |(datain[307:304] ^ 12);
  assign w796[2] = |(datain[303:300] ^ 3);
  assign w796[3] = |(datain[299:296] ^ 5);
  assign w796[4] = |(datain[295:292] ^ 12);
  assign w796[5] = |(datain[291:288] ^ 13);
  assign w796[6] = |(datain[287:284] ^ 2);
  assign w796[7] = |(datain[283:280] ^ 1);
  assign w796[8] = |(datain[279:276] ^ 2);
  assign w796[9] = |(datain[275:272] ^ 6);
  assign w796[10] = |(datain[271:268] ^ 8);
  assign w796[11] = |(datain[267:264] ^ 11);
  assign w796[12] = |(datain[263:260] ^ 4);
  assign w796[13] = |(datain[259:256] ^ 7);
  assign w796[14] = |(datain[255:252] ^ 15);
  assign w796[15] = |(datain[251:248] ^ 14);
  assign w796[16] = |(datain[247:244] ^ 2);
  assign w796[17] = |(datain[243:240] ^ 14);
  assign w796[18] = |(datain[239:236] ^ 3);
  assign w796[19] = |(datain[235:232] ^ 11);
  assign w796[20] = |(datain[231:228] ^ 0);
  assign w796[21] = |(datain[227:224] ^ 6);
  assign w796[22] = |(datain[223:220] ^ 14);
  assign w796[23] = |(datain[219:216] ^ 14);
  assign w796[24] = |(datain[215:212] ^ 0);
  assign w796[25] = |(datain[211:208] ^ 2);
  assign w796[26] = |(datain[207:204] ^ 7);
  assign w796[27] = |(datain[203:200] ^ 4);
  assign w796[28] = |(datain[199:196] ^ 3);
  assign w796[29] = |(datain[195:192] ^ 1);
  assign w796[30] = |(datain[191:188] ^ 8);
  assign w796[31] = |(datain[187:184] ^ 9);
  assign comp[796] = ~(|w796);
  wire [28-1:0] w797;
  assign w797[0] = |(datain[311:308] ^ 13);
  assign w797[1] = |(datain[307:304] ^ 3);
  assign w797[2] = |(datain[303:300] ^ 14);
  assign w797[3] = |(datain[299:296] ^ 11);
  assign w797[4] = |(datain[295:292] ^ 2);
  assign w797[5] = |(datain[291:288] ^ 4);
  assign w797[6] = |(datain[287:284] ^ 0);
  assign w797[7] = |(datain[283:280] ^ 15);
  assign w797[8] = |(datain[279:276] ^ 3);
  assign w797[9] = |(datain[275:272] ^ 12);
  assign w797[10] = |(datain[271:268] ^ 0);
  assign w797[11] = |(datain[267:264] ^ 0);
  assign w797[12] = |(datain[263:260] ^ 7);
  assign w797[13] = |(datain[259:256] ^ 4);
  assign w797[14] = |(datain[255:252] ^ 0);
  assign w797[15] = |(datain[251:248] ^ 1);
  assign w797[16] = |(datain[247:244] ^ 4);
  assign w797[17] = |(datain[243:240] ^ 3);
  assign w797[18] = |(datain[239:236] ^ 8);
  assign w797[19] = |(datain[235:232] ^ 9);
  assign w797[20] = |(datain[231:228] ^ 1);
  assign w797[21] = |(datain[227:224] ^ 14);
  assign w797[22] = |(datain[223:220] ^ 0);
  assign w797[23] = |(datain[219:216] ^ 12);
  assign w797[24] = |(datain[215:212] ^ 0);
  assign w797[25] = |(datain[211:208] ^ 0);
  assign w797[26] = |(datain[207:204] ^ 12);
  assign w797[27] = |(datain[203:200] ^ 7);
  assign comp[797] = ~(|w797);
  wire [40-1:0] w798;
  assign w798[0] = |(datain[311:308] ^ 4);
  assign w798[1] = |(datain[307:304] ^ 2);
  assign w798[2] = |(datain[303:300] ^ 3);
  assign w798[3] = |(datain[299:296] ^ 3);
  assign w798[4] = |(datain[295:292] ^ 12);
  assign w798[5] = |(datain[291:288] ^ 9);
  assign w798[6] = |(datain[287:284] ^ 3);
  assign w798[7] = |(datain[283:280] ^ 3);
  assign w798[8] = |(datain[279:276] ^ 13);
  assign w798[9] = |(datain[275:272] ^ 2);
  assign w798[10] = |(datain[271:268] ^ 8);
  assign w798[11] = |(datain[267:264] ^ 11);
  assign w798[12] = |(datain[263:260] ^ 1);
  assign w798[13] = |(datain[259:256] ^ 14);
  assign w798[14] = |(datain[255:252] ^ 1);
  assign w798[15] = |(datain[251:248] ^ 12);
  assign w798[16] = |(datain[247:244] ^ 0);
  assign w798[17] = |(datain[243:240] ^ 0);
  assign w798[18] = |(datain[239:236] ^ 12);
  assign w798[19] = |(datain[235:232] ^ 13);
  assign w798[20] = |(datain[231:228] ^ 2);
  assign w798[21] = |(datain[227:224] ^ 1);
  assign w798[22] = |(datain[223:220] ^ 11);
  assign w798[23] = |(datain[219:216] ^ 4);
  assign w798[24] = |(datain[215:212] ^ 4);
  assign w798[25] = |(datain[211:208] ^ 0);
  assign w798[26] = |(datain[207:204] ^ 8);
  assign w798[27] = |(datain[203:200] ^ 13);
  assign w798[28] = |(datain[199:196] ^ 1);
  assign w798[29] = |(datain[195:192] ^ 6);
  assign w798[30] = |(datain[191:188] ^ 0);
  assign w798[31] = |(datain[187:184] ^ 0);
  assign w798[32] = |(datain[183:180] ^ 0);
  assign w798[33] = |(datain[179:176] ^ 0);
  assign w798[34] = |(datain[175:172] ^ 11);
  assign w798[35] = |(datain[171:168] ^ 9);
  assign w798[36] = |(datain[167:164] ^ 0);
  assign w798[37] = |(datain[163:160] ^ 14);
  assign w798[38] = |(datain[159:156] ^ 0);
  assign w798[39] = |(datain[155:152] ^ 0);
  assign comp[798] = ~(|w798);
  wire [48-1:0] w799;
  assign w799[0] = |(datain[311:308] ^ 11);
  assign w799[1] = |(datain[307:304] ^ 15);
  assign w799[2] = |(datain[303:300] ^ 0);
  assign w799[3] = |(datain[299:296] ^ 0);
  assign w799[4] = |(datain[295:292] ^ 0);
  assign w799[5] = |(datain[291:288] ^ 1);
  assign w799[6] = |(datain[287:284] ^ 15);
  assign w799[7] = |(datain[283:280] ^ 3);
  assign w799[8] = |(datain[279:276] ^ 10);
  assign w799[9] = |(datain[275:272] ^ 4);
  assign w799[10] = |(datain[271:268] ^ 11);
  assign w799[11] = |(datain[267:264] ^ 8);
  assign w799[12] = |(datain[263:260] ^ 13);
  assign w799[13] = |(datain[259:256] ^ 10);
  assign w799[14] = |(datain[255:252] ^ 11);
  assign w799[15] = |(datain[251:248] ^ 14);
  assign w799[16] = |(datain[247:244] ^ 12);
  assign w799[17] = |(datain[243:240] ^ 13);
  assign w799[18] = |(datain[239:236] ^ 2);
  assign w799[19] = |(datain[235:232] ^ 1);
  assign w799[20] = |(datain[231:228] ^ 3);
  assign w799[21] = |(datain[227:224] ^ 13);
  assign w799[22] = |(datain[223:220] ^ 15);
  assign w799[23] = |(datain[219:216] ^ 14);
  assign w799[24] = |(datain[215:212] ^ 12);
  assign w799[25] = |(datain[211:208] ^ 0);
  assign w799[26] = |(datain[207:204] ^ 7);
  assign w799[27] = |(datain[203:200] ^ 5);
  assign w799[28] = |(datain[199:196] ^ 0);
  assign w799[29] = |(datain[195:192] ^ 3);
  assign w799[30] = |(datain[191:188] ^ 14);
  assign w799[31] = |(datain[187:184] ^ 11);
  assign w799[32] = |(datain[183:180] ^ 7);
  assign w799[33] = |(datain[179:176] ^ 3);
  assign w799[34] = |(datain[175:172] ^ 9);
  assign w799[35] = |(datain[171:168] ^ 0);
  assign w799[36] = |(datain[167:164] ^ 11);
  assign w799[37] = |(datain[163:160] ^ 4);
  assign w799[38] = |(datain[159:156] ^ 5);
  assign w799[39] = |(datain[155:152] ^ 2);
  assign w799[40] = |(datain[151:148] ^ 12);
  assign w799[41] = |(datain[147:144] ^ 13);
  assign w799[42] = |(datain[143:140] ^ 2);
  assign w799[43] = |(datain[139:136] ^ 1);
  assign w799[44] = |(datain[135:132] ^ 2);
  assign w799[45] = |(datain[131:128] ^ 6);
  assign w799[46] = |(datain[127:124] ^ 8);
  assign w799[47] = |(datain[123:120] ^ 11);
  assign comp[799] = ~(|w799);
  wire [74-1:0] w800;
  assign w800[0] = |(datain[311:308] ^ 14);
  assign w800[1] = |(datain[307:304] ^ 11);
  assign w800[2] = |(datain[303:300] ^ 0);
  assign w800[3] = |(datain[299:296] ^ 6);
  assign w800[4] = |(datain[295:292] ^ 11);
  assign w800[5] = |(datain[291:288] ^ 9);
  assign w800[6] = |(datain[287:284] ^ 1);
  assign w800[7] = |(datain[283:280] ^ 8);
  assign w800[8] = |(datain[279:276] ^ 0);
  assign w800[9] = |(datain[275:272] ^ 0);
  assign w800[10] = |(datain[271:268] ^ 12);
  assign w800[11] = |(datain[267:264] ^ 13);
  assign w800[12] = |(datain[263:260] ^ 2);
  assign w800[13] = |(datain[259:256] ^ 1);
  assign w800[14] = |(datain[255:252] ^ 14);
  assign w800[15] = |(datain[251:248] ^ 11);
  assign w800[16] = |(datain[247:244] ^ 1);
  assign w800[17] = |(datain[243:240] ^ 3);
  assign w800[18] = |(datain[239:236] ^ 11);
  assign w800[19] = |(datain[235:232] ^ 8);
  assign w800[20] = |(datain[231:228] ^ 0);
  assign w800[21] = |(datain[227:224] ^ 2);
  assign w800[22] = |(datain[223:220] ^ 4);
  assign w800[23] = |(datain[219:216] ^ 2);
  assign w800[24] = |(datain[215:212] ^ 3);
  assign w800[25] = |(datain[211:208] ^ 3);
  assign w800[26] = |(datain[207:204] ^ 12);
  assign w800[27] = |(datain[203:200] ^ 9);
  assign w800[28] = |(datain[199:196] ^ 3);
  assign w800[29] = |(datain[195:192] ^ 3);
  assign w800[30] = |(datain[191:188] ^ 13);
  assign w800[31] = |(datain[187:184] ^ 2);
  assign w800[32] = |(datain[183:180] ^ 12);
  assign w800[33] = |(datain[179:176] ^ 13);
  assign w800[34] = |(datain[175:172] ^ 2);
  assign w800[35] = |(datain[171:168] ^ 1);
  assign w800[36] = |(datain[167:164] ^ 11);
  assign w800[37] = |(datain[163:160] ^ 9);
  assign w800[38] = |(datain[159:156] ^ 15);
  assign w800[39] = |(datain[155:152] ^ 10);
  assign w800[40] = |(datain[151:148] ^ 0);
  assign w800[41] = |(datain[147:144] ^ 5);
  assign w800[42] = |(datain[143:140] ^ 9);
  assign w800[43] = |(datain[139:136] ^ 0);
  assign w800[44] = |(datain[135:132] ^ 11);
  assign w800[45] = |(datain[131:128] ^ 10);
  assign w800[46] = |(datain[127:124] ^ 1);
  assign w800[47] = |(datain[123:120] ^ 0);
  assign w800[48] = |(datain[119:116] ^ 0);
  assign w800[49] = |(datain[115:112] ^ 1);
  assign w800[50] = |(datain[111:108] ^ 14);
  assign w800[51] = |(datain[107:104] ^ 8);
  assign w800[52] = |(datain[103:100] ^ 2);
  assign w800[53] = |(datain[99:96] ^ 11);
  assign w800[54] = |(datain[95:92] ^ 0);
  assign w800[55] = |(datain[91:88] ^ 1);
  assign w800[56] = |(datain[87:84] ^ 11);
  assign w800[57] = |(datain[83:80] ^ 8);
  assign w800[58] = |(datain[79:76] ^ 0);
  assign w800[59] = |(datain[75:72] ^ 1);
  assign w800[60] = |(datain[71:68] ^ 5);
  assign w800[61] = |(datain[67:64] ^ 7);
  assign w800[62] = |(datain[63:60] ^ 11);
  assign w800[63] = |(datain[59:56] ^ 9);
  assign w800[64] = |(datain[55:52] ^ 13);
  assign w800[65] = |(datain[51:48] ^ 10);
  assign w800[66] = |(datain[47:44] ^ 11);
  assign w800[67] = |(datain[43:40] ^ 14);
  assign w800[68] = |(datain[39:36] ^ 8);
  assign w800[69] = |(datain[35:32] ^ 11);
  assign w800[70] = |(datain[31:28] ^ 1);
  assign w800[71] = |(datain[27:24] ^ 6);
  assign w800[72] = |(datain[23:20] ^ 11);
  assign w800[73] = |(datain[19:16] ^ 9);
  assign comp[800] = ~(|w800);
  wire [42-1:0] w801;
  assign w801[0] = |(datain[311:308] ^ 15);
  assign w801[1] = |(datain[307:304] ^ 3);
  assign w801[2] = |(datain[303:300] ^ 10);
  assign w801[3] = |(datain[299:296] ^ 4);
  assign w801[4] = |(datain[295:292] ^ 11);
  assign w801[5] = |(datain[291:288] ^ 8);
  assign w801[6] = |(datain[287:284] ^ 13);
  assign w801[7] = |(datain[283:280] ^ 10);
  assign w801[8] = |(datain[279:276] ^ 11);
  assign w801[9] = |(datain[275:272] ^ 14);
  assign w801[10] = |(datain[271:268] ^ 12);
  assign w801[11] = |(datain[267:264] ^ 13);
  assign w801[12] = |(datain[263:260] ^ 2);
  assign w801[13] = |(datain[259:256] ^ 1);
  assign w801[14] = |(datain[255:252] ^ 3);
  assign w801[15] = |(datain[251:248] ^ 13);
  assign w801[16] = |(datain[247:244] ^ 15);
  assign w801[17] = |(datain[243:240] ^ 14);
  assign w801[18] = |(datain[239:236] ^ 12);
  assign w801[19] = |(datain[235:232] ^ 0);
  assign w801[20] = |(datain[231:228] ^ 7);
  assign w801[21] = |(datain[227:224] ^ 5);
  assign w801[22] = |(datain[223:220] ^ 0);
  assign w801[23] = |(datain[219:216] ^ 3);
  assign w801[24] = |(datain[215:212] ^ 14);
  assign w801[25] = |(datain[211:208] ^ 11);
  assign w801[26] = |(datain[207:204] ^ 5);
  assign w801[27] = |(datain[203:200] ^ 14);
  assign w801[28] = |(datain[199:196] ^ 9);
  assign w801[29] = |(datain[195:192] ^ 0);
  assign w801[30] = |(datain[191:188] ^ 11);
  assign w801[31] = |(datain[187:184] ^ 4);
  assign w801[32] = |(datain[183:180] ^ 5);
  assign w801[33] = |(datain[179:176] ^ 2);
  assign w801[34] = |(datain[175:172] ^ 12);
  assign w801[35] = |(datain[171:168] ^ 13);
  assign w801[36] = |(datain[167:164] ^ 2);
  assign w801[37] = |(datain[163:160] ^ 1);
  assign w801[38] = |(datain[159:156] ^ 2);
  assign w801[39] = |(datain[155:152] ^ 6);
  assign w801[40] = |(datain[151:148] ^ 8);
  assign w801[41] = |(datain[147:144] ^ 11);
  assign comp[801] = ~(|w801);
  wire [46-1:0] w802;
  assign w802[0] = |(datain[311:308] ^ 4);
  assign w802[1] = |(datain[307:304] ^ 0);
  assign w802[2] = |(datain[303:300] ^ 14);
  assign w802[3] = |(datain[299:296] ^ 11);
  assign w802[4] = |(datain[295:292] ^ 0);
  assign w802[5] = |(datain[291:288] ^ 2);
  assign w802[6] = |(datain[287:284] ^ 11);
  assign w802[7] = |(datain[283:280] ^ 4);
  assign w802[8] = |(datain[279:276] ^ 3);
  assign w802[9] = |(datain[275:272] ^ 15);
  assign w802[10] = |(datain[271:268] ^ 14);
  assign w802[11] = |(datain[267:264] ^ 8);
  assign w802[12] = |(datain[263:260] ^ 1);
  assign w802[13] = |(datain[259:256] ^ 5);
  assign w802[14] = |(datain[255:252] ^ 0);
  assign w802[15] = |(datain[251:248] ^ 0);
  assign w802[16] = |(datain[247:244] ^ 7);
  assign w802[17] = |(datain[243:240] ^ 2);
  assign w802[18] = |(datain[239:236] ^ 0);
  assign w802[19] = |(datain[235:232] ^ 2);
  assign w802[20] = |(datain[231:228] ^ 2);
  assign w802[21] = |(datain[227:224] ^ 11);
  assign w802[22] = |(datain[223:220] ^ 12);
  assign w802[23] = |(datain[219:216] ^ 1);
  assign w802[24] = |(datain[215:212] ^ 12);
  assign w802[25] = |(datain[211:208] ^ 3);
  assign w802[26] = |(datain[207:204] ^ 3);
  assign w802[27] = |(datain[203:200] ^ 3);
  assign w802[28] = |(datain[199:196] ^ 12);
  assign w802[29] = |(datain[195:192] ^ 9);
  assign w802[30] = |(datain[191:188] ^ 3);
  assign w802[31] = |(datain[187:184] ^ 3);
  assign w802[32] = |(datain[183:180] ^ 13);
  assign w802[33] = |(datain[179:176] ^ 2);
  assign w802[34] = |(datain[175:172] ^ 11);
  assign w802[35] = |(datain[171:168] ^ 8);
  assign w802[36] = |(datain[167:164] ^ 0);
  assign w802[37] = |(datain[163:160] ^ 2);
  assign w802[38] = |(datain[159:156] ^ 4);
  assign w802[39] = |(datain[155:152] ^ 2);
  assign w802[40] = |(datain[151:148] ^ 14);
  assign w802[41] = |(datain[147:144] ^ 11);
  assign w802[42] = |(datain[143:140] ^ 0);
  assign w802[43] = |(datain[139:136] ^ 7);
  assign w802[44] = |(datain[135:132] ^ 3);
  assign w802[45] = |(datain[131:128] ^ 3);
  assign comp[802] = ~(|w802);
  wire [74-1:0] w803;
  assign w803[0] = |(datain[311:308] ^ 10);
  assign w803[1] = |(datain[307:304] ^ 11);
  assign w803[2] = |(datain[303:300] ^ 5);
  assign w803[3] = |(datain[299:296] ^ 8);
  assign w803[4] = |(datain[295:292] ^ 2);
  assign w803[5] = |(datain[291:288] ^ 13);
  assign w803[6] = |(datain[287:284] ^ 0);
  assign w803[7] = |(datain[283:280] ^ 4);
  assign w803[8] = |(datain[279:276] ^ 0);
  assign w803[9] = |(datain[275:272] ^ 0);
  assign w803[10] = |(datain[271:268] ^ 10);
  assign w803[11] = |(datain[267:264] ^ 11);
  assign w803[12] = |(datain[263:260] ^ 11);
  assign w803[13] = |(datain[259:256] ^ 4);
  assign w803[14] = |(datain[255:252] ^ 4);
  assign w803[15] = |(datain[251:248] ^ 0);
  assign w803[16] = |(datain[247:244] ^ 11);
  assign w803[17] = |(datain[243:240] ^ 9);
  assign w803[18] = |(datain[239:236] ^ 1);
  assign w803[19] = |(datain[235:232] ^ 0);
  assign w803[20] = |(datain[231:228] ^ 0);
  assign w803[21] = |(datain[227:224] ^ 1);
  assign w803[22] = |(datain[223:220] ^ 3);
  assign w803[23] = |(datain[219:216] ^ 3);
  assign w803[24] = |(datain[215:212] ^ 13);
  assign w803[25] = |(datain[211:208] ^ 2);
  assign w803[26] = |(datain[207:204] ^ 12);
  assign w803[27] = |(datain[203:200] ^ 13);
  assign w803[28] = |(datain[199:196] ^ 2);
  assign w803[29] = |(datain[195:192] ^ 1);
  assign w803[30] = |(datain[191:188] ^ 3);
  assign w803[31] = |(datain[187:184] ^ 2);
  assign w803[32] = |(datain[183:180] ^ 12);
  assign w803[33] = |(datain[179:176] ^ 0);
  assign w803[34] = |(datain[175:172] ^ 14);
  assign w803[35] = |(datain[171:168] ^ 8);
  assign w803[36] = |(datain[167:164] ^ 6);
  assign w803[37] = |(datain[163:160] ^ 4);
  assign w803[38] = |(datain[159:156] ^ 15);
  assign w803[39] = |(datain[155:152] ^ 15);
  assign w803[40] = |(datain[151:148] ^ 11);
  assign w803[41] = |(datain[147:144] ^ 4);
  assign w803[42] = |(datain[143:140] ^ 4);
  assign w803[43] = |(datain[139:136] ^ 0);
  assign w803[44] = |(datain[135:132] ^ 11);
  assign w803[45] = |(datain[131:128] ^ 9);
  assign w803[46] = |(datain[127:124] ^ 1);
  assign w803[47] = |(datain[123:120] ^ 8);
  assign w803[48] = |(datain[119:116] ^ 0);
  assign w803[49] = |(datain[115:112] ^ 0);
  assign w803[50] = |(datain[111:108] ^ 11);
  assign w803[51] = |(datain[107:104] ^ 10);
  assign w803[52] = |(datain[103:100] ^ 1);
  assign w803[53] = |(datain[99:96] ^ 4);
  assign w803[54] = |(datain[95:92] ^ 0);
  assign w803[55] = |(datain[91:88] ^ 1);
  assign w803[56] = |(datain[87:84] ^ 12);
  assign w803[57] = |(datain[83:80] ^ 13);
  assign w803[58] = |(datain[79:76] ^ 2);
  assign w803[59] = |(datain[75:72] ^ 1);
  assign w803[60] = |(datain[71:68] ^ 11);
  assign w803[61] = |(datain[67:64] ^ 4);
  assign w803[62] = |(datain[63:60] ^ 3);
  assign w803[63] = |(datain[59:56] ^ 14);
  assign w803[64] = |(datain[55:52] ^ 12);
  assign w803[65] = |(datain[51:48] ^ 13);
  assign w803[66] = |(datain[47:44] ^ 2);
  assign w803[67] = |(datain[43:40] ^ 1);
  assign w803[68] = |(datain[39:36] ^ 0);
  assign w803[69] = |(datain[35:32] ^ 7);
  assign w803[70] = |(datain[31:28] ^ 1);
  assign w803[71] = |(datain[27:24] ^ 15);
  assign w803[72] = |(datain[23:20] ^ 6);
  assign w803[73] = |(datain[19:16] ^ 1);
  assign comp[803] = ~(|w803);
  wire [76-1:0] w804;
  assign w804[0] = |(datain[311:308] ^ 11);
  assign w804[1] = |(datain[307:304] ^ 9);
  assign w804[2] = |(datain[303:300] ^ 11);
  assign w804[3] = |(datain[299:296] ^ 7);
  assign w804[4] = |(datain[295:292] ^ 0);
  assign w804[5] = |(datain[291:288] ^ 1);
  assign w804[6] = |(datain[287:284] ^ 11);
  assign w804[7] = |(datain[283:280] ^ 4);
  assign w804[8] = |(datain[279:276] ^ 4);
  assign w804[9] = |(datain[275:272] ^ 0);
  assign w804[10] = |(datain[271:268] ^ 14);
  assign w804[11] = |(datain[267:264] ^ 8);
  assign w804[12] = |(datain[263:260] ^ 13);
  assign w804[13] = |(datain[259:256] ^ 10);
  assign w804[14] = |(datain[255:252] ^ 0);
  assign w804[15] = |(datain[251:248] ^ 0);
  assign w804[16] = |(datain[247:244] ^ 3);
  assign w804[17] = |(datain[243:240] ^ 9);
  assign w804[18] = |(datain[239:236] ^ 12);
  assign w804[19] = |(datain[235:232] ^ 8);
  assign w804[20] = |(datain[231:228] ^ 7);
  assign w804[21] = |(datain[227:224] ^ 5);
  assign w804[22] = |(datain[223:220] ^ 0);
  assign w804[23] = |(datain[219:216] ^ 14);
  assign w804[24] = |(datain[215:212] ^ 14);
  assign w804[25] = |(datain[211:208] ^ 8);
  assign w804[26] = |(datain[207:204] ^ 4);
  assign w804[27] = |(datain[203:200] ^ 8);
  assign w804[28] = |(datain[199:196] ^ 0);
  assign w804[29] = |(datain[195:192] ^ 0);
  assign w804[30] = |(datain[191:188] ^ 11);
  assign w804[31] = |(datain[187:184] ^ 10);
  assign w804[32] = |(datain[183:180] ^ 11);
  assign w804[33] = |(datain[179:176] ^ 4);
  assign w804[34] = |(datain[175:172] ^ 0);
  assign w804[35] = |(datain[171:168] ^ 1);
  assign w804[36] = |(datain[167:164] ^ 11);
  assign w804[37] = |(datain[163:160] ^ 9);
  assign w804[38] = |(datain[159:156] ^ 0);
  assign w804[39] = |(datain[155:152] ^ 3);
  assign w804[40] = |(datain[151:148] ^ 0);
  assign w804[41] = |(datain[147:144] ^ 0);
  assign w804[42] = |(datain[143:140] ^ 11);
  assign w804[43] = |(datain[139:136] ^ 4);
  assign w804[44] = |(datain[135:132] ^ 4);
  assign w804[45] = |(datain[131:128] ^ 0);
  assign w804[46] = |(datain[127:124] ^ 14);
  assign w804[47] = |(datain[123:120] ^ 8);
  assign w804[48] = |(datain[119:116] ^ 12);
  assign w804[49] = |(datain[115:112] ^ 8);
  assign w804[50] = |(datain[111:108] ^ 0);
  assign w804[51] = |(datain[107:104] ^ 0);
  assign w804[52] = |(datain[103:100] ^ 11);
  assign w804[53] = |(datain[99:96] ^ 8);
  assign w804[54] = |(datain[95:92] ^ 0);
  assign w804[55] = |(datain[91:88] ^ 1);
  assign w804[56] = |(datain[87:84] ^ 5);
  assign w804[57] = |(datain[83:80] ^ 7);
  assign w804[58] = |(datain[79:76] ^ 8);
  assign w804[59] = |(datain[75:72] ^ 11);
  assign w804[60] = |(datain[71:68] ^ 0);
  assign w804[61] = |(datain[67:64] ^ 14);
  assign w804[62] = |(datain[63:60] ^ 11);
  assign w804[63] = |(datain[59:56] ^ 10);
  assign w804[64] = |(datain[55:52] ^ 0);
  assign w804[65] = |(datain[51:48] ^ 1);
  assign w804[66] = |(datain[47:44] ^ 8);
  assign w804[67] = |(datain[43:40] ^ 11);
  assign w804[68] = |(datain[39:36] ^ 1);
  assign w804[69] = |(datain[35:32] ^ 6);
  assign w804[70] = |(datain[31:28] ^ 11);
  assign w804[71] = |(datain[27:24] ^ 12);
  assign w804[72] = |(datain[23:20] ^ 0);
  assign w804[73] = |(datain[19:16] ^ 1);
  assign w804[74] = |(datain[15:12] ^ 14);
  assign w804[75] = |(datain[11:8] ^ 8);
  assign comp[804] = ~(|w804);
  wire [48-1:0] w805;
  assign w805[0] = |(datain[311:308] ^ 5);
  assign w805[1] = |(datain[307:304] ^ 0);
  assign w805[2] = |(datain[303:300] ^ 2);
  assign w805[3] = |(datain[299:296] ^ 13);
  assign w805[4] = |(datain[295:292] ^ 0);
  assign w805[5] = |(datain[291:288] ^ 0);
  assign w805[6] = |(datain[287:284] ^ 4);
  assign w805[7] = |(datain[283:280] ^ 11);
  assign w805[8] = |(datain[279:276] ^ 7);
  assign w805[9] = |(datain[275:272] ^ 4);
  assign w805[10] = |(datain[271:268] ^ 7);
  assign w805[11] = |(datain[267:264] ^ 6);
  assign w805[12] = |(datain[263:260] ^ 5);
  assign w805[13] = |(datain[259:256] ^ 8);
  assign w805[14] = |(datain[255:252] ^ 5);
  assign w805[15] = |(datain[251:248] ^ 0);
  assign w805[16] = |(datain[247:244] ^ 8);
  assign w805[17] = |(datain[243:240] ^ 0);
  assign w805[18] = |(datain[239:236] ^ 14);
  assign w805[19] = |(datain[235:232] ^ 12);
  assign w805[20] = |(datain[231:228] ^ 4);
  assign w805[21] = |(datain[227:224] ^ 14);
  assign w805[22] = |(datain[223:220] ^ 7);
  assign w805[23] = |(datain[219:216] ^ 4);
  assign w805[24] = |(datain[215:212] ^ 0);
  assign w805[25] = |(datain[211:208] ^ 10);
  assign w805[26] = |(datain[207:204] ^ 5);
  assign w805[27] = |(datain[203:200] ^ 8);
  assign w805[28] = |(datain[199:196] ^ 5);
  assign w805[29] = |(datain[195:192] ^ 0);
  assign w805[30] = |(datain[191:188] ^ 8);
  assign w805[31] = |(datain[187:184] ^ 0);
  assign w805[32] = |(datain[183:180] ^ 14);
  assign w805[33] = |(datain[179:176] ^ 12);
  assign w805[34] = |(datain[175:172] ^ 4);
  assign w805[35] = |(datain[171:168] ^ 15);
  assign w805[36] = |(datain[167:164] ^ 7);
  assign w805[37] = |(datain[163:160] ^ 4);
  assign w805[38] = |(datain[159:156] ^ 0);
  assign w805[39] = |(datain[155:152] ^ 3);
  assign w805[40] = |(datain[151:148] ^ 14);
  assign w805[41] = |(datain[147:144] ^ 9);
  assign w805[42] = |(datain[143:140] ^ 8);
  assign w805[43] = |(datain[139:136] ^ 11);
  assign w805[44] = |(datain[135:132] ^ 0);
  assign w805[45] = |(datain[131:128] ^ 2);
  assign w805[46] = |(datain[127:124] ^ 2);
  assign w805[47] = |(datain[123:120] ^ 14);
  assign comp[805] = ~(|w805);
  wire [76-1:0] w806;
  assign w806[0] = |(datain[311:308] ^ 0);
  assign w806[1] = |(datain[307:304] ^ 3);
  assign w806[2] = |(datain[303:300] ^ 11);
  assign w806[3] = |(datain[299:296] ^ 9);
  assign w806[4] = |(datain[295:292] ^ 10);
  assign w806[5] = |(datain[291:288] ^ 12);
  assign w806[6] = |(datain[287:284] ^ 0);
  assign w806[7] = |(datain[283:280] ^ 10);
  assign w806[8] = |(datain[279:276] ^ 2);
  assign w806[9] = |(datain[275:272] ^ 11);
  assign w806[10] = |(datain[271:268] ^ 12);
  assign w806[11] = |(datain[267:264] ^ 11);
  assign w806[12] = |(datain[263:260] ^ 2);
  assign w806[13] = |(datain[259:256] ^ 14);
  assign w806[14] = |(datain[255:252] ^ 10);
  assign w806[15] = |(datain[251:248] ^ 0);
  assign w806[16] = |(datain[247:244] ^ 13);
  assign w806[17] = |(datain[243:240] ^ 14);
  assign w806[18] = |(datain[239:236] ^ 0);
  assign w806[19] = |(datain[235:232] ^ 1);
  assign w806[20] = |(datain[231:228] ^ 2);
  assign w806[21] = |(datain[227:224] ^ 14);
  assign w806[22] = |(datain[223:220] ^ 3);
  assign w806[23] = |(datain[219:216] ^ 0);
  assign w806[24] = |(datain[215:212] ^ 0);
  assign w806[25] = |(datain[211:208] ^ 7);
  assign w806[26] = |(datain[207:204] ^ 4);
  assign w806[27] = |(datain[203:200] ^ 3);
  assign w806[28] = |(datain[199:196] ^ 14);
  assign w806[29] = |(datain[195:192] ^ 2);
  assign w806[30] = |(datain[191:188] ^ 15);
  assign w806[31] = |(datain[187:184] ^ 10);
  assign w806[32] = |(datain[183:180] ^ 9);
  assign w806[33] = |(datain[179:176] ^ 13);
  assign w806[34] = |(datain[175:172] ^ 5);
  assign w806[35] = |(datain[171:168] ^ 8);
  assign w806[36] = |(datain[167:164] ^ 5);
  assign w806[37] = |(datain[163:160] ^ 9);
  assign w806[38] = |(datain[159:156] ^ 5);
  assign w806[39] = |(datain[155:152] ^ 11);
  assign w806[40] = |(datain[151:148] ^ 12);
  assign w806[41] = |(datain[147:144] ^ 3);
  assign w806[42] = |(datain[143:140] ^ 14);
  assign w806[43] = |(datain[139:136] ^ 8);
  assign w806[44] = |(datain[135:132] ^ 14);
  assign w806[45] = |(datain[131:128] ^ 2);
  assign w806[46] = |(datain[127:124] ^ 15);
  assign w806[47] = |(datain[123:120] ^ 15);
  assign w806[48] = |(datain[119:116] ^ 11);
  assign w806[49] = |(datain[115:112] ^ 4);
  assign w806[50] = |(datain[111:108] ^ 4);
  assign w806[51] = |(datain[107:104] ^ 0);
  assign w806[52] = |(datain[103:100] ^ 11);
  assign w806[53] = |(datain[99:96] ^ 9);
  assign w806[54] = |(datain[95:92] ^ 10);
  assign w806[55] = |(datain[91:88] ^ 12);
  assign w806[56] = |(datain[87:84] ^ 0);
  assign w806[57] = |(datain[83:80] ^ 10);
  assign w806[58] = |(datain[79:76] ^ 11);
  assign w806[59] = |(datain[75:72] ^ 10);
  assign w806[60] = |(datain[71:68] ^ 0);
  assign w806[61] = |(datain[67:64] ^ 3);
  assign w806[62] = |(datain[63:60] ^ 0);
  assign w806[63] = |(datain[59:56] ^ 1);
  assign w806[64] = |(datain[55:52] ^ 2);
  assign w806[65] = |(datain[51:48] ^ 11);
  assign w806[66] = |(datain[47:44] ^ 12);
  assign w806[67] = |(datain[43:40] ^ 10);
  assign w806[68] = |(datain[39:36] ^ 8);
  assign w806[69] = |(datain[35:32] ^ 11);
  assign w806[70] = |(datain[31:28] ^ 1);
  assign w806[71] = |(datain[27:24] ^ 14);
  assign w806[72] = |(datain[23:20] ^ 12);
  assign w806[73] = |(datain[19:16] ^ 4);
  assign w806[74] = |(datain[15:12] ^ 0);
  assign w806[75] = |(datain[11:8] ^ 10);
  assign comp[806] = ~(|w806);
  wire [76-1:0] w807;
  assign w807[0] = |(datain[311:308] ^ 0);
  assign w807[1] = |(datain[307:304] ^ 2);
  assign w807[2] = |(datain[303:300] ^ 11);
  assign w807[3] = |(datain[299:296] ^ 9);
  assign w807[4] = |(datain[295:292] ^ 3);
  assign w807[5] = |(datain[291:288] ^ 15);
  assign w807[6] = |(datain[287:284] ^ 0);
  assign w807[7] = |(datain[283:280] ^ 11);
  assign w807[8] = |(datain[279:276] ^ 2);
  assign w807[9] = |(datain[275:272] ^ 11);
  assign w807[10] = |(datain[271:268] ^ 12);
  assign w807[11] = |(datain[267:264] ^ 11);
  assign w807[12] = |(datain[263:260] ^ 2);
  assign w807[13] = |(datain[259:256] ^ 14);
  assign w807[14] = |(datain[255:252] ^ 10);
  assign w807[15] = |(datain[251:248] ^ 0);
  assign w807[16] = |(datain[247:244] ^ 13);
  assign w807[17] = |(datain[243:240] ^ 14);
  assign w807[18] = |(datain[239:236] ^ 0);
  assign w807[19] = |(datain[235:232] ^ 1);
  assign w807[20] = |(datain[231:228] ^ 2);
  assign w807[21] = |(datain[227:224] ^ 14);
  assign w807[22] = |(datain[223:220] ^ 3);
  assign w807[23] = |(datain[219:216] ^ 0);
  assign w807[24] = |(datain[215:212] ^ 0);
  assign w807[25] = |(datain[211:208] ^ 7);
  assign w807[26] = |(datain[207:204] ^ 4);
  assign w807[27] = |(datain[203:200] ^ 3);
  assign w807[28] = |(datain[199:196] ^ 14);
  assign w807[29] = |(datain[195:192] ^ 2);
  assign w807[30] = |(datain[191:188] ^ 15);
  assign w807[31] = |(datain[187:184] ^ 10);
  assign w807[32] = |(datain[183:180] ^ 9);
  assign w807[33] = |(datain[179:176] ^ 13);
  assign w807[34] = |(datain[175:172] ^ 5);
  assign w807[35] = |(datain[171:168] ^ 8);
  assign w807[36] = |(datain[167:164] ^ 5);
  assign w807[37] = |(datain[163:160] ^ 9);
  assign w807[38] = |(datain[159:156] ^ 5);
  assign w807[39] = |(datain[155:152] ^ 11);
  assign w807[40] = |(datain[151:148] ^ 12);
  assign w807[41] = |(datain[147:144] ^ 3);
  assign w807[42] = |(datain[143:140] ^ 14);
  assign w807[43] = |(datain[139:136] ^ 8);
  assign w807[44] = |(datain[135:132] ^ 14);
  assign w807[45] = |(datain[131:128] ^ 2);
  assign w807[46] = |(datain[127:124] ^ 15);
  assign w807[47] = |(datain[123:120] ^ 15);
  assign w807[48] = |(datain[119:116] ^ 11);
  assign w807[49] = |(datain[115:112] ^ 4);
  assign w807[50] = |(datain[111:108] ^ 4);
  assign w807[51] = |(datain[107:104] ^ 0);
  assign w807[52] = |(datain[103:100] ^ 11);
  assign w807[53] = |(datain[99:96] ^ 9);
  assign w807[54] = |(datain[95:92] ^ 3);
  assign w807[55] = |(datain[91:88] ^ 15);
  assign w807[56] = |(datain[87:84] ^ 0);
  assign w807[57] = |(datain[83:80] ^ 11);
  assign w807[58] = |(datain[79:76] ^ 11);
  assign w807[59] = |(datain[75:72] ^ 10);
  assign w807[60] = |(datain[71:68] ^ 0);
  assign w807[61] = |(datain[67:64] ^ 3);
  assign w807[62] = |(datain[63:60] ^ 0);
  assign w807[63] = |(datain[59:56] ^ 1);
  assign w807[64] = |(datain[55:52] ^ 2);
  assign w807[65] = |(datain[51:48] ^ 11);
  assign w807[66] = |(datain[47:44] ^ 12);
  assign w807[67] = |(datain[43:40] ^ 10);
  assign w807[68] = |(datain[39:36] ^ 8);
  assign w807[69] = |(datain[35:32] ^ 11);
  assign w807[70] = |(datain[31:28] ^ 1);
  assign w807[71] = |(datain[27:24] ^ 14);
  assign w807[72] = |(datain[23:20] ^ 5);
  assign w807[73] = |(datain[19:16] ^ 8);
  assign w807[74] = |(datain[15:12] ^ 0);
  assign w807[75] = |(datain[11:8] ^ 11);
  assign comp[807] = ~(|w807);
  wire [76-1:0] w808;
  assign w808[0] = |(datain[311:308] ^ 0);
  assign w808[1] = |(datain[307:304] ^ 12);
  assign w808[2] = |(datain[303:300] ^ 2);
  assign w808[3] = |(datain[299:296] ^ 11);
  assign w808[4] = |(datain[295:292] ^ 12);
  assign w808[5] = |(datain[291:288] ^ 11);
  assign w808[6] = |(datain[287:284] ^ 2);
  assign w808[7] = |(datain[283:280] ^ 14);
  assign w808[8] = |(datain[279:276] ^ 10);
  assign w808[9] = |(datain[275:272] ^ 0);
  assign w808[10] = |(datain[271:268] ^ 13);
  assign w808[11] = |(datain[267:264] ^ 14);
  assign w808[12] = |(datain[263:260] ^ 0);
  assign w808[13] = |(datain[259:256] ^ 1);
  assign w808[14] = |(datain[255:252] ^ 2);
  assign w808[15] = |(datain[251:248] ^ 14);
  assign w808[16] = |(datain[247:244] ^ 3);
  assign w808[17] = |(datain[243:240] ^ 0);
  assign w808[18] = |(datain[239:236] ^ 0);
  assign w808[19] = |(datain[235:232] ^ 7);
  assign w808[20] = |(datain[231:228] ^ 4);
  assign w808[21] = |(datain[227:224] ^ 3);
  assign w808[22] = |(datain[223:220] ^ 14);
  assign w808[23] = |(datain[219:216] ^ 2);
  assign w808[24] = |(datain[215:212] ^ 15);
  assign w808[25] = |(datain[211:208] ^ 10);
  assign w808[26] = |(datain[207:204] ^ 9);
  assign w808[27] = |(datain[203:200] ^ 13);
  assign w808[28] = |(datain[199:196] ^ 5);
  assign w808[29] = |(datain[195:192] ^ 8);
  assign w808[30] = |(datain[191:188] ^ 5);
  assign w808[31] = |(datain[187:184] ^ 9);
  assign w808[32] = |(datain[183:180] ^ 5);
  assign w808[33] = |(datain[179:176] ^ 11);
  assign w808[34] = |(datain[175:172] ^ 12);
  assign w808[35] = |(datain[171:168] ^ 3);
  assign w808[36] = |(datain[167:164] ^ 14);
  assign w808[37] = |(datain[163:160] ^ 8);
  assign w808[38] = |(datain[159:156] ^ 14);
  assign w808[39] = |(datain[155:152] ^ 2);
  assign w808[40] = |(datain[151:148] ^ 15);
  assign w808[41] = |(datain[147:144] ^ 15);
  assign w808[42] = |(datain[143:140] ^ 11);
  assign w808[43] = |(datain[139:136] ^ 4);
  assign w808[44] = |(datain[135:132] ^ 4);
  assign w808[45] = |(datain[131:128] ^ 0);
  assign w808[46] = |(datain[127:124] ^ 11);
  assign w808[47] = |(datain[123:120] ^ 9);
  assign w808[48] = |(datain[119:116] ^ 2);
  assign w808[49] = |(datain[115:112] ^ 5);
  assign w808[50] = |(datain[111:108] ^ 0);
  assign w808[51] = |(datain[107:104] ^ 12);
  assign w808[52] = |(datain[103:100] ^ 11);
  assign w808[53] = |(datain[99:96] ^ 10);
  assign w808[54] = |(datain[95:92] ^ 0);
  assign w808[55] = |(datain[91:88] ^ 3);
  assign w808[56] = |(datain[87:84] ^ 0);
  assign w808[57] = |(datain[83:80] ^ 1);
  assign w808[58] = |(datain[79:76] ^ 2);
  assign w808[59] = |(datain[75:72] ^ 11);
  assign w808[60] = |(datain[71:68] ^ 12);
  assign w808[61] = |(datain[67:64] ^ 10);
  assign w808[62] = |(datain[63:60] ^ 8);
  assign w808[63] = |(datain[59:56] ^ 11);
  assign w808[64] = |(datain[55:52] ^ 1);
  assign w808[65] = |(datain[51:48] ^ 14);
  assign w808[66] = |(datain[47:44] ^ 3);
  assign w808[67] = |(datain[43:40] ^ 14);
  assign w808[68] = |(datain[39:36] ^ 0);
  assign w808[69] = |(datain[35:32] ^ 12);
  assign w808[70] = |(datain[31:28] ^ 14);
  assign w808[71] = |(datain[27:24] ^ 8);
  assign w808[72] = |(datain[23:20] ^ 6);
  assign w808[73] = |(datain[19:16] ^ 0);
  assign w808[74] = |(datain[15:12] ^ 0);
  assign w808[75] = |(datain[11:8] ^ 0);
  assign comp[808] = ~(|w808);
  wire [66-1:0] w809;
  assign w809[0] = |(datain[311:308] ^ 15);
  assign w809[1] = |(datain[307:304] ^ 10);
  assign w809[2] = |(datain[303:300] ^ 9);
  assign w809[3] = |(datain[299:296] ^ 13);
  assign w809[4] = |(datain[295:292] ^ 5);
  assign w809[5] = |(datain[291:288] ^ 8);
  assign w809[6] = |(datain[287:284] ^ 5);
  assign w809[7] = |(datain[283:280] ^ 9);
  assign w809[8] = |(datain[279:276] ^ 5);
  assign w809[9] = |(datain[275:272] ^ 11);
  assign w809[10] = |(datain[271:268] ^ 12);
  assign w809[11] = |(datain[267:264] ^ 3);
  assign w809[12] = |(datain[263:260] ^ 14);
  assign w809[13] = |(datain[259:256] ^ 8);
  assign w809[14] = |(datain[255:252] ^ 14);
  assign w809[15] = |(datain[251:248] ^ 2);
  assign w809[16] = |(datain[247:244] ^ 15);
  assign w809[17] = |(datain[243:240] ^ 15);
  assign w809[18] = |(datain[239:236] ^ 11);
  assign w809[19] = |(datain[235:232] ^ 4);
  assign w809[20] = |(datain[231:228] ^ 4);
  assign w809[21] = |(datain[227:224] ^ 0);
  assign w809[22] = |(datain[223:220] ^ 11);
  assign w809[23] = |(datain[219:216] ^ 9);
  assign w809[24] = |(datain[215:212] ^ 9);
  assign w809[25] = |(datain[211:208] ^ 9);
  assign w809[26] = |(datain[207:204] ^ 0);
  assign w809[27] = |(datain[203:200] ^ 12);
  assign w809[28] = |(datain[199:196] ^ 11);
  assign w809[29] = |(datain[195:192] ^ 10);
  assign w809[30] = |(datain[191:188] ^ 0);
  assign w809[31] = |(datain[187:184] ^ 3);
  assign w809[32] = |(datain[183:180] ^ 0);
  assign w809[33] = |(datain[179:176] ^ 1);
  assign w809[34] = |(datain[175:172] ^ 2);
  assign w809[35] = |(datain[171:168] ^ 11);
  assign w809[36] = |(datain[167:164] ^ 12);
  assign w809[37] = |(datain[163:160] ^ 10);
  assign w809[38] = |(datain[159:156] ^ 8);
  assign w809[39] = |(datain[155:152] ^ 11);
  assign w809[40] = |(datain[151:148] ^ 1);
  assign w809[41] = |(datain[147:144] ^ 14);
  assign w809[42] = |(datain[143:140] ^ 11);
  assign w809[43] = |(datain[139:136] ^ 2);
  assign w809[44] = |(datain[135:132] ^ 0);
  assign w809[45] = |(datain[131:128] ^ 12);
  assign w809[46] = |(datain[127:124] ^ 14);
  assign w809[47] = |(datain[123:120] ^ 8);
  assign w809[48] = |(datain[119:116] ^ 14);
  assign w809[49] = |(datain[115:112] ^ 15);
  assign w809[50] = |(datain[111:108] ^ 0);
  assign w809[51] = |(datain[107:104] ^ 0);
  assign w809[52] = |(datain[103:100] ^ 14);
  assign w809[53] = |(datain[99:96] ^ 8);
  assign w809[54] = |(datain[95:92] ^ 12);
  assign w809[55] = |(datain[91:88] ^ 14);
  assign w809[56] = |(datain[87:84] ^ 15);
  assign w809[57] = |(datain[83:80] ^ 15);
  assign w809[58] = |(datain[79:76] ^ 12);
  assign w809[59] = |(datain[75:72] ^ 3);
  assign w809[60] = |(datain[71:68] ^ 11);
  assign w809[61] = |(datain[67:64] ^ 0);
  assign w809[62] = |(datain[63:60] ^ 0);
  assign w809[63] = |(datain[59:56] ^ 3);
  assign w809[64] = |(datain[55:52] ^ 12);
  assign w809[65] = |(datain[51:48] ^ 15);
  assign comp[809] = ~(|w809);
  wire [46-1:0] w810;
  assign w810[0] = |(datain[311:308] ^ 9);
  assign w810[1] = |(datain[307:304] ^ 0);
  assign w810[2] = |(datain[303:300] ^ 8);
  assign w810[3] = |(datain[299:296] ^ 0);
  assign w810[4] = |(datain[295:292] ^ 15);
  assign w810[5] = |(datain[291:288] ^ 12);
  assign w810[6] = |(datain[287:284] ^ 3);
  assign w810[7] = |(datain[283:280] ^ 11);
  assign w810[8] = |(datain[279:276] ^ 7);
  assign w810[9] = |(datain[275:272] ^ 5);
  assign w810[10] = |(datain[271:268] ^ 0);
  assign w810[11] = |(datain[267:264] ^ 3);
  assign w810[12] = |(datain[263:260] ^ 14);
  assign w810[13] = |(datain[259:256] ^ 9);
  assign w810[14] = |(datain[255:252] ^ 7);
  assign w810[15] = |(datain[251:248] ^ 2);
  assign w810[16] = |(datain[247:244] ^ 15);
  assign w810[17] = |(datain[243:240] ^ 15);
  assign w810[18] = |(datain[239:236] ^ 3);
  assign w810[19] = |(datain[235:232] ^ 13);
  assign w810[20] = |(datain[231:228] ^ 0);
  assign w810[21] = |(datain[227:224] ^ 0);
  assign w810[22] = |(datain[223:220] ^ 3);
  assign w810[23] = |(datain[219:216] ^ 13);
  assign w810[24] = |(datain[215:212] ^ 7);
  assign w810[25] = |(datain[211:208] ^ 4);
  assign w810[26] = |(datain[207:204] ^ 0);
  assign w810[27] = |(datain[203:200] ^ 15);
  assign w810[28] = |(datain[199:196] ^ 3);
  assign w810[29] = |(datain[195:192] ^ 13);
  assign w810[30] = |(datain[191:188] ^ 0);
  assign w810[31] = |(datain[187:184] ^ 2);
  assign w810[32] = |(datain[183:180] ^ 3);
  assign w810[33] = |(datain[179:176] ^ 13);
  assign w810[34] = |(datain[175:172] ^ 7);
  assign w810[35] = |(datain[171:168] ^ 4);
  assign w810[36] = |(datain[167:164] ^ 0);
  assign w810[37] = |(datain[163:160] ^ 10);
  assign w810[38] = |(datain[159:156] ^ 8);
  assign w810[39] = |(datain[155:152] ^ 0);
  assign w810[40] = |(datain[151:148] ^ 15);
  assign w810[41] = |(datain[147:144] ^ 12);
  assign w810[42] = |(datain[143:140] ^ 5);
  assign w810[43] = |(datain[139:136] ^ 6);
  assign w810[44] = |(datain[135:132] ^ 7);
  assign w810[45] = |(datain[131:128] ^ 4);
  assign comp[810] = ~(|w810);
  wire [72-1:0] w811;
  assign w811[0] = |(datain[311:308] ^ 12);
  assign w811[1] = |(datain[307:304] ^ 11);
  assign w811[2] = |(datain[303:300] ^ 2);
  assign w811[3] = |(datain[299:296] ^ 14);
  assign w811[4] = |(datain[295:292] ^ 10);
  assign w811[5] = |(datain[291:288] ^ 0);
  assign w811[6] = |(datain[287:284] ^ 13);
  assign w811[7] = |(datain[283:280] ^ 2);
  assign w811[8] = |(datain[279:276] ^ 0);
  assign w811[9] = |(datain[275:272] ^ 1);
  assign w811[10] = |(datain[271:268] ^ 2);
  assign w811[11] = |(datain[267:264] ^ 14);
  assign w811[12] = |(datain[263:260] ^ 3);
  assign w811[13] = |(datain[259:256] ^ 0);
  assign w811[14] = |(datain[255:252] ^ 0);
  assign w811[15] = |(datain[251:248] ^ 7);
  assign w811[16] = |(datain[247:244] ^ 4);
  assign w811[17] = |(datain[243:240] ^ 3);
  assign w811[18] = |(datain[239:236] ^ 14);
  assign w811[19] = |(datain[235:232] ^ 2);
  assign w811[20] = |(datain[231:228] ^ 15);
  assign w811[21] = |(datain[227:224] ^ 10);
  assign w811[22] = |(datain[223:220] ^ 9);
  assign w811[23] = |(datain[219:216] ^ 13);
  assign w811[24] = |(datain[215:212] ^ 5);
  assign w811[25] = |(datain[211:208] ^ 8);
  assign w811[26] = |(datain[207:204] ^ 5);
  assign w811[27] = |(datain[203:200] ^ 9);
  assign w811[28] = |(datain[199:196] ^ 5);
  assign w811[29] = |(datain[195:192] ^ 11);
  assign w811[30] = |(datain[191:188] ^ 12);
  assign w811[31] = |(datain[187:184] ^ 3);
  assign w811[32] = |(datain[183:180] ^ 14);
  assign w811[33] = |(datain[179:176] ^ 8);
  assign w811[34] = |(datain[175:172] ^ 14);
  assign w811[35] = |(datain[171:168] ^ 2);
  assign w811[36] = |(datain[167:164] ^ 15);
  assign w811[37] = |(datain[163:160] ^ 15);
  assign w811[38] = |(datain[159:156] ^ 11);
  assign w811[39] = |(datain[155:152] ^ 4);
  assign w811[40] = |(datain[151:148] ^ 4);
  assign w811[41] = |(datain[147:144] ^ 0);
  assign w811[42] = |(datain[143:140] ^ 11);
  assign w811[43] = |(datain[139:136] ^ 9);
  assign w811[44] = |(datain[135:132] ^ 2);
  assign w811[45] = |(datain[131:128] ^ 3);
  assign w811[46] = |(datain[127:124] ^ 0);
  assign w811[47] = |(datain[123:120] ^ 14);
  assign w811[48] = |(datain[119:116] ^ 11);
  assign w811[49] = |(datain[115:112] ^ 10);
  assign w811[50] = |(datain[111:108] ^ 0);
  assign w811[51] = |(datain[107:104] ^ 3);
  assign w811[52] = |(datain[103:100] ^ 0);
  assign w811[53] = |(datain[99:96] ^ 1);
  assign w811[54] = |(datain[95:92] ^ 2);
  assign w811[55] = |(datain[91:88] ^ 11);
  assign w811[56] = |(datain[87:84] ^ 12);
  assign w811[57] = |(datain[83:80] ^ 10);
  assign w811[58] = |(datain[79:76] ^ 8);
  assign w811[59] = |(datain[75:72] ^ 11);
  assign w811[60] = |(datain[71:68] ^ 1);
  assign w811[61] = |(datain[67:64] ^ 14);
  assign w811[62] = |(datain[63:60] ^ 3);
  assign w811[63] = |(datain[59:56] ^ 12);
  assign w811[64] = |(datain[55:52] ^ 0);
  assign w811[65] = |(datain[51:48] ^ 14);
  assign w811[66] = |(datain[47:44] ^ 14);
  assign w811[67] = |(datain[43:40] ^ 8);
  assign w811[68] = |(datain[39:36] ^ 2);
  assign w811[69] = |(datain[35:32] ^ 4);
  assign w811[70] = |(datain[31:28] ^ 0);
  assign w811[71] = |(datain[27:24] ^ 1);
  assign comp[811] = ~(|w811);
  wire [72-1:0] w812;
  assign w812[0] = |(datain[311:308] ^ 12);
  assign w812[1] = |(datain[307:304] ^ 11);
  assign w812[2] = |(datain[303:300] ^ 2);
  assign w812[3] = |(datain[299:296] ^ 14);
  assign w812[4] = |(datain[295:292] ^ 10);
  assign w812[5] = |(datain[291:288] ^ 0);
  assign w812[6] = |(datain[287:284] ^ 13);
  assign w812[7] = |(datain[283:280] ^ 13);
  assign w812[8] = |(datain[279:276] ^ 0);
  assign w812[9] = |(datain[275:272] ^ 1);
  assign w812[10] = |(datain[271:268] ^ 2);
  assign w812[11] = |(datain[267:264] ^ 14);
  assign w812[12] = |(datain[263:260] ^ 3);
  assign w812[13] = |(datain[259:256] ^ 0);
  assign w812[14] = |(datain[255:252] ^ 0);
  assign w812[15] = |(datain[251:248] ^ 7);
  assign w812[16] = |(datain[247:244] ^ 4);
  assign w812[17] = |(datain[243:240] ^ 3);
  assign w812[18] = |(datain[239:236] ^ 14);
  assign w812[19] = |(datain[235:232] ^ 2);
  assign w812[20] = |(datain[231:228] ^ 15);
  assign w812[21] = |(datain[227:224] ^ 10);
  assign w812[22] = |(datain[223:220] ^ 9);
  assign w812[23] = |(datain[219:216] ^ 13);
  assign w812[24] = |(datain[215:212] ^ 5);
  assign w812[25] = |(datain[211:208] ^ 8);
  assign w812[26] = |(datain[207:204] ^ 5);
  assign w812[27] = |(datain[203:200] ^ 9);
  assign w812[28] = |(datain[199:196] ^ 5);
  assign w812[29] = |(datain[195:192] ^ 11);
  assign w812[30] = |(datain[191:188] ^ 12);
  assign w812[31] = |(datain[187:184] ^ 3);
  assign w812[32] = |(datain[183:180] ^ 14);
  assign w812[33] = |(datain[179:176] ^ 8);
  assign w812[34] = |(datain[175:172] ^ 14);
  assign w812[35] = |(datain[171:168] ^ 2);
  assign w812[36] = |(datain[167:164] ^ 15);
  assign w812[37] = |(datain[163:160] ^ 15);
  assign w812[38] = |(datain[159:156] ^ 11);
  assign w812[39] = |(datain[155:152] ^ 4);
  assign w812[40] = |(datain[151:148] ^ 4);
  assign w812[41] = |(datain[147:144] ^ 0);
  assign w812[42] = |(datain[143:140] ^ 11);
  assign w812[43] = |(datain[139:136] ^ 9);
  assign w812[44] = |(datain[135:132] ^ 12);
  assign w812[45] = |(datain[131:128] ^ 5);
  assign w812[46] = |(datain[127:124] ^ 0);
  assign w812[47] = |(datain[123:120] ^ 14);
  assign w812[48] = |(datain[119:116] ^ 11);
  assign w812[49] = |(datain[115:112] ^ 10);
  assign w812[50] = |(datain[111:108] ^ 0);
  assign w812[51] = |(datain[107:104] ^ 3);
  assign w812[52] = |(datain[103:100] ^ 0);
  assign w812[53] = |(datain[99:96] ^ 1);
  assign w812[54] = |(datain[95:92] ^ 2);
  assign w812[55] = |(datain[91:88] ^ 11);
  assign w812[56] = |(datain[87:84] ^ 12);
  assign w812[57] = |(datain[83:80] ^ 10);
  assign w812[58] = |(datain[79:76] ^ 8);
  assign w812[59] = |(datain[75:72] ^ 11);
  assign w812[60] = |(datain[71:68] ^ 1);
  assign w812[61] = |(datain[67:64] ^ 14);
  assign w812[62] = |(datain[63:60] ^ 13);
  assign w812[63] = |(datain[59:56] ^ 14);
  assign w812[64] = |(datain[55:52] ^ 0);
  assign w812[65] = |(datain[51:48] ^ 14);
  assign w812[66] = |(datain[47:44] ^ 14);
  assign w812[67] = |(datain[43:40] ^ 8);
  assign w812[68] = |(datain[39:36] ^ 13);
  assign w812[69] = |(datain[35:32] ^ 2);
  assign w812[70] = |(datain[31:28] ^ 0);
  assign w812[71] = |(datain[27:24] ^ 1);
  assign comp[812] = ~(|w812);
  wire [72-1:0] w813;
  assign w813[0] = |(datain[311:308] ^ 12);
  assign w813[1] = |(datain[307:304] ^ 11);
  assign w813[2] = |(datain[303:300] ^ 2);
  assign w813[3] = |(datain[299:296] ^ 14);
  assign w813[4] = |(datain[295:292] ^ 10);
  assign w813[5] = |(datain[291:288] ^ 0);
  assign w813[6] = |(datain[287:284] ^ 13);
  assign w813[7] = |(datain[283:280] ^ 13);
  assign w813[8] = |(datain[279:276] ^ 0);
  assign w813[9] = |(datain[275:272] ^ 1);
  assign w813[10] = |(datain[271:268] ^ 2);
  assign w813[11] = |(datain[267:264] ^ 14);
  assign w813[12] = |(datain[263:260] ^ 3);
  assign w813[13] = |(datain[259:256] ^ 0);
  assign w813[14] = |(datain[255:252] ^ 0);
  assign w813[15] = |(datain[251:248] ^ 7);
  assign w813[16] = |(datain[247:244] ^ 4);
  assign w813[17] = |(datain[243:240] ^ 3);
  assign w813[18] = |(datain[239:236] ^ 14);
  assign w813[19] = |(datain[235:232] ^ 2);
  assign w813[20] = |(datain[231:228] ^ 15);
  assign w813[21] = |(datain[227:224] ^ 10);
  assign w813[22] = |(datain[223:220] ^ 9);
  assign w813[23] = |(datain[219:216] ^ 13);
  assign w813[24] = |(datain[215:212] ^ 5);
  assign w813[25] = |(datain[211:208] ^ 8);
  assign w813[26] = |(datain[207:204] ^ 5);
  assign w813[27] = |(datain[203:200] ^ 9);
  assign w813[28] = |(datain[199:196] ^ 5);
  assign w813[29] = |(datain[195:192] ^ 11);
  assign w813[30] = |(datain[191:188] ^ 12);
  assign w813[31] = |(datain[187:184] ^ 3);
  assign w813[32] = |(datain[183:180] ^ 14);
  assign w813[33] = |(datain[179:176] ^ 8);
  assign w813[34] = |(datain[175:172] ^ 14);
  assign w813[35] = |(datain[171:168] ^ 2);
  assign w813[36] = |(datain[167:164] ^ 15);
  assign w813[37] = |(datain[163:160] ^ 15);
  assign w813[38] = |(datain[159:156] ^ 11);
  assign w813[39] = |(datain[155:152] ^ 4);
  assign w813[40] = |(datain[151:148] ^ 4);
  assign w813[41] = |(datain[147:144] ^ 0);
  assign w813[42] = |(datain[143:140] ^ 11);
  assign w813[43] = |(datain[139:136] ^ 9);
  assign w813[44] = |(datain[135:132] ^ 1);
  assign w813[45] = |(datain[131:128] ^ 15);
  assign w813[46] = |(datain[127:124] ^ 0);
  assign w813[47] = |(datain[123:120] ^ 15);
  assign w813[48] = |(datain[119:116] ^ 11);
  assign w813[49] = |(datain[115:112] ^ 10);
  assign w813[50] = |(datain[111:108] ^ 0);
  assign w813[51] = |(datain[107:104] ^ 3);
  assign w813[52] = |(datain[103:100] ^ 0);
  assign w813[53] = |(datain[99:96] ^ 1);
  assign w813[54] = |(datain[95:92] ^ 2);
  assign w813[55] = |(datain[91:88] ^ 11);
  assign w813[56] = |(datain[87:84] ^ 12);
  assign w813[57] = |(datain[83:80] ^ 10);
  assign w813[58] = |(datain[79:76] ^ 8);
  assign w813[59] = |(datain[75:72] ^ 11);
  assign w813[60] = |(datain[71:68] ^ 1);
  assign w813[61] = |(datain[67:64] ^ 14);
  assign w813[62] = |(datain[63:60] ^ 3);
  assign w813[63] = |(datain[59:56] ^ 8);
  assign w813[64] = |(datain[55:52] ^ 0);
  assign w813[65] = |(datain[51:48] ^ 15);
  assign w813[66] = |(datain[47:44] ^ 14);
  assign w813[67] = |(datain[43:40] ^ 8);
  assign w813[68] = |(datain[39:36] ^ 4);
  assign w813[69] = |(datain[35:32] ^ 6);
  assign w813[70] = |(datain[31:28] ^ 0);
  assign w813[71] = |(datain[27:24] ^ 1);
  assign comp[813] = ~(|w813);
  wire [74-1:0] w814;
  assign w814[0] = |(datain[311:308] ^ 11);
  assign w814[1] = |(datain[307:304] ^ 9);
  assign w814[2] = |(datain[303:300] ^ 5);
  assign w814[3] = |(datain[299:296] ^ 15);
  assign w814[4] = |(datain[295:292] ^ 0);
  assign w814[5] = |(datain[291:288] ^ 13);
  assign w814[6] = |(datain[287:284] ^ 2);
  assign w814[7] = |(datain[283:280] ^ 11);
  assign w814[8] = |(datain[279:276] ^ 12);
  assign w814[9] = |(datain[275:272] ^ 11);
  assign w814[10] = |(datain[271:268] ^ 2);
  assign w814[11] = |(datain[267:264] ^ 14);
  assign w814[12] = |(datain[263:260] ^ 10);
  assign w814[13] = |(datain[259:256] ^ 0);
  assign w814[14] = |(datain[255:252] ^ 13);
  assign w814[15] = |(datain[251:248] ^ 14);
  assign w814[16] = |(datain[247:244] ^ 0);
  assign w814[17] = |(datain[243:240] ^ 1);
  assign w814[18] = |(datain[239:236] ^ 2);
  assign w814[19] = |(datain[235:232] ^ 14);
  assign w814[20] = |(datain[231:228] ^ 3);
  assign w814[21] = |(datain[227:224] ^ 0);
  assign w814[22] = |(datain[223:220] ^ 0);
  assign w814[23] = |(datain[219:216] ^ 7);
  assign w814[24] = |(datain[215:212] ^ 4);
  assign w814[25] = |(datain[211:208] ^ 3);
  assign w814[26] = |(datain[207:204] ^ 14);
  assign w814[27] = |(datain[203:200] ^ 2);
  assign w814[28] = |(datain[199:196] ^ 15);
  assign w814[29] = |(datain[195:192] ^ 10);
  assign w814[30] = |(datain[191:188] ^ 9);
  assign w814[31] = |(datain[187:184] ^ 13);
  assign w814[32] = |(datain[183:180] ^ 5);
  assign w814[33] = |(datain[179:176] ^ 8);
  assign w814[34] = |(datain[175:172] ^ 5);
  assign w814[35] = |(datain[171:168] ^ 9);
  assign w814[36] = |(datain[167:164] ^ 5);
  assign w814[37] = |(datain[163:160] ^ 11);
  assign w814[38] = |(datain[159:156] ^ 12);
  assign w814[39] = |(datain[155:152] ^ 3);
  assign w814[40] = |(datain[151:148] ^ 14);
  assign w814[41] = |(datain[147:144] ^ 8);
  assign w814[42] = |(datain[143:140] ^ 14);
  assign w814[43] = |(datain[139:136] ^ 2);
  assign w814[44] = |(datain[135:132] ^ 15);
  assign w814[45] = |(datain[131:128] ^ 15);
  assign w814[46] = |(datain[127:124] ^ 11);
  assign w814[47] = |(datain[123:120] ^ 4);
  assign w814[48] = |(datain[119:116] ^ 4);
  assign w814[49] = |(datain[115:112] ^ 0);
  assign w814[50] = |(datain[111:108] ^ 11);
  assign w814[51] = |(datain[107:104] ^ 9);
  assign w814[52] = |(datain[103:100] ^ 5);
  assign w814[53] = |(datain[99:96] ^ 15);
  assign w814[54] = |(datain[95:92] ^ 0);
  assign w814[55] = |(datain[91:88] ^ 13);
  assign w814[56] = |(datain[87:84] ^ 11);
  assign w814[57] = |(datain[83:80] ^ 10);
  assign w814[58] = |(datain[79:76] ^ 0);
  assign w814[59] = |(datain[75:72] ^ 3);
  assign w814[60] = |(datain[71:68] ^ 0);
  assign w814[61] = |(datain[67:64] ^ 1);
  assign w814[62] = |(datain[63:60] ^ 2);
  assign w814[63] = |(datain[59:56] ^ 11);
  assign w814[64] = |(datain[55:52] ^ 12);
  assign w814[65] = |(datain[51:48] ^ 10);
  assign w814[66] = |(datain[47:44] ^ 8);
  assign w814[67] = |(datain[43:40] ^ 11);
  assign w814[68] = |(datain[39:36] ^ 1);
  assign w814[69] = |(datain[35:32] ^ 14);
  assign w814[70] = |(datain[31:28] ^ 7);
  assign w814[71] = |(datain[27:24] ^ 8);
  assign w814[72] = |(datain[23:20] ^ 0);
  assign w814[73] = |(datain[19:16] ^ 13);
  assign comp[814] = ~(|w814);
  wire [46-1:0] w815;
  assign w815[0] = |(datain[311:308] ^ 9);
  assign w815[1] = |(datain[307:304] ^ 0);
  assign w815[2] = |(datain[303:300] ^ 8);
  assign w815[3] = |(datain[299:296] ^ 0);
  assign w815[4] = |(datain[295:292] ^ 15);
  assign w815[5] = |(datain[291:288] ^ 12);
  assign w815[6] = |(datain[287:284] ^ 3);
  assign w815[7] = |(datain[283:280] ^ 11);
  assign w815[8] = |(datain[279:276] ^ 7);
  assign w815[9] = |(datain[275:272] ^ 5);
  assign w815[10] = |(datain[271:268] ^ 0);
  assign w815[11] = |(datain[267:264] ^ 3);
  assign w815[12] = |(datain[263:260] ^ 14);
  assign w815[13] = |(datain[259:256] ^ 9);
  assign w815[14] = |(datain[255:252] ^ 1);
  assign w815[15] = |(datain[251:248] ^ 8);
  assign w815[16] = |(datain[247:244] ^ 15);
  assign w815[17] = |(datain[243:240] ^ 15);
  assign w815[18] = |(datain[239:236] ^ 3);
  assign w815[19] = |(datain[235:232] ^ 13);
  assign w815[20] = |(datain[231:228] ^ 0);
  assign w815[21] = |(datain[227:224] ^ 0);
  assign w815[22] = |(datain[223:220] ^ 3);
  assign w815[23] = |(datain[219:216] ^ 13);
  assign w815[24] = |(datain[215:212] ^ 7);
  assign w815[25] = |(datain[211:208] ^ 4);
  assign w815[26] = |(datain[207:204] ^ 0);
  assign w815[27] = |(datain[203:200] ^ 15);
  assign w815[28] = |(datain[199:196] ^ 3);
  assign w815[29] = |(datain[195:192] ^ 13);
  assign w815[30] = |(datain[191:188] ^ 0);
  assign w815[31] = |(datain[187:184] ^ 2);
  assign w815[32] = |(datain[183:180] ^ 3);
  assign w815[33] = |(datain[179:176] ^ 13);
  assign w815[34] = |(datain[175:172] ^ 7);
  assign w815[35] = |(datain[171:168] ^ 4);
  assign w815[36] = |(datain[167:164] ^ 0);
  assign w815[37] = |(datain[163:160] ^ 10);
  assign w815[38] = |(datain[159:156] ^ 8);
  assign w815[39] = |(datain[155:152] ^ 0);
  assign w815[40] = |(datain[151:148] ^ 15);
  assign w815[41] = |(datain[147:144] ^ 12);
  assign w815[42] = |(datain[143:140] ^ 5);
  assign w815[43] = |(datain[139:136] ^ 6);
  assign w815[44] = |(datain[135:132] ^ 7);
  assign w815[45] = |(datain[131:128] ^ 4);
  assign comp[815] = ~(|w815);
  wire [74-1:0] w816;
  assign w816[0] = |(datain[311:308] ^ 11);
  assign w816[1] = |(datain[307:304] ^ 9);
  assign w816[2] = |(datain[303:300] ^ 7);
  assign w816[3] = |(datain[299:296] ^ 11);
  assign w816[4] = |(datain[295:292] ^ 0);
  assign w816[5] = |(datain[291:288] ^ 13);
  assign w816[6] = |(datain[287:284] ^ 2);
  assign w816[7] = |(datain[283:280] ^ 11);
  assign w816[8] = |(datain[279:276] ^ 12);
  assign w816[9] = |(datain[275:272] ^ 11);
  assign w816[10] = |(datain[271:268] ^ 2);
  assign w816[11] = |(datain[267:264] ^ 14);
  assign w816[12] = |(datain[263:260] ^ 10);
  assign w816[13] = |(datain[259:256] ^ 0);
  assign w816[14] = |(datain[255:252] ^ 13);
  assign w816[15] = |(datain[251:248] ^ 14);
  assign w816[16] = |(datain[247:244] ^ 0);
  assign w816[17] = |(datain[243:240] ^ 1);
  assign w816[18] = |(datain[239:236] ^ 2);
  assign w816[19] = |(datain[235:232] ^ 14);
  assign w816[20] = |(datain[231:228] ^ 3);
  assign w816[21] = |(datain[227:224] ^ 0);
  assign w816[22] = |(datain[223:220] ^ 0);
  assign w816[23] = |(datain[219:216] ^ 7);
  assign w816[24] = |(datain[215:212] ^ 4);
  assign w816[25] = |(datain[211:208] ^ 3);
  assign w816[26] = |(datain[207:204] ^ 14);
  assign w816[27] = |(datain[203:200] ^ 2);
  assign w816[28] = |(datain[199:196] ^ 15);
  assign w816[29] = |(datain[195:192] ^ 10);
  assign w816[30] = |(datain[191:188] ^ 9);
  assign w816[31] = |(datain[187:184] ^ 13);
  assign w816[32] = |(datain[183:180] ^ 5);
  assign w816[33] = |(datain[179:176] ^ 8);
  assign w816[34] = |(datain[175:172] ^ 5);
  assign w816[35] = |(datain[171:168] ^ 9);
  assign w816[36] = |(datain[167:164] ^ 5);
  assign w816[37] = |(datain[163:160] ^ 11);
  assign w816[38] = |(datain[159:156] ^ 12);
  assign w816[39] = |(datain[155:152] ^ 3);
  assign w816[40] = |(datain[151:148] ^ 14);
  assign w816[41] = |(datain[147:144] ^ 8);
  assign w816[42] = |(datain[143:140] ^ 14);
  assign w816[43] = |(datain[139:136] ^ 2);
  assign w816[44] = |(datain[135:132] ^ 15);
  assign w816[45] = |(datain[131:128] ^ 15);
  assign w816[46] = |(datain[127:124] ^ 11);
  assign w816[47] = |(datain[123:120] ^ 4);
  assign w816[48] = |(datain[119:116] ^ 4);
  assign w816[49] = |(datain[115:112] ^ 0);
  assign w816[50] = |(datain[111:108] ^ 11);
  assign w816[51] = |(datain[107:104] ^ 9);
  assign w816[52] = |(datain[103:100] ^ 7);
  assign w816[53] = |(datain[99:96] ^ 11);
  assign w816[54] = |(datain[95:92] ^ 0);
  assign w816[55] = |(datain[91:88] ^ 13);
  assign w816[56] = |(datain[87:84] ^ 11);
  assign w816[57] = |(datain[83:80] ^ 10);
  assign w816[58] = |(datain[79:76] ^ 0);
  assign w816[59] = |(datain[75:72] ^ 3);
  assign w816[60] = |(datain[71:68] ^ 0);
  assign w816[61] = |(datain[67:64] ^ 1);
  assign w816[62] = |(datain[63:60] ^ 2);
  assign w816[63] = |(datain[59:56] ^ 11);
  assign w816[64] = |(datain[55:52] ^ 12);
  assign w816[65] = |(datain[51:48] ^ 10);
  assign w816[66] = |(datain[47:44] ^ 8);
  assign w816[67] = |(datain[43:40] ^ 11);
  assign w816[68] = |(datain[39:36] ^ 1);
  assign w816[69] = |(datain[35:32] ^ 14);
  assign w816[70] = |(datain[31:28] ^ 9);
  assign w816[71] = |(datain[27:24] ^ 4);
  assign w816[72] = |(datain[23:20] ^ 0);
  assign w816[73] = |(datain[19:16] ^ 13);
  assign comp[816] = ~(|w816);
  wire [72-1:0] w817;
  assign w817[0] = |(datain[311:308] ^ 12);
  assign w817[1] = |(datain[307:304] ^ 11);
  assign w817[2] = |(datain[303:300] ^ 2);
  assign w817[3] = |(datain[299:296] ^ 14);
  assign w817[4] = |(datain[295:292] ^ 10);
  assign w817[5] = |(datain[291:288] ^ 0);
  assign w817[6] = |(datain[287:284] ^ 13);
  assign w817[7] = |(datain[283:280] ^ 12);
  assign w817[8] = |(datain[279:276] ^ 0);
  assign w817[9] = |(datain[275:272] ^ 1);
  assign w817[10] = |(datain[271:268] ^ 2);
  assign w817[11] = |(datain[267:264] ^ 14);
  assign w817[12] = |(datain[263:260] ^ 3);
  assign w817[13] = |(datain[259:256] ^ 0);
  assign w817[14] = |(datain[255:252] ^ 0);
  assign w817[15] = |(datain[251:248] ^ 7);
  assign w817[16] = |(datain[247:244] ^ 4);
  assign w817[17] = |(datain[243:240] ^ 3);
  assign w817[18] = |(datain[239:236] ^ 14);
  assign w817[19] = |(datain[235:232] ^ 2);
  assign w817[20] = |(datain[231:228] ^ 15);
  assign w817[21] = |(datain[227:224] ^ 10);
  assign w817[22] = |(datain[223:220] ^ 9);
  assign w817[23] = |(datain[219:216] ^ 13);
  assign w817[24] = |(datain[215:212] ^ 5);
  assign w817[25] = |(datain[211:208] ^ 8);
  assign w817[26] = |(datain[207:204] ^ 5);
  assign w817[27] = |(datain[203:200] ^ 9);
  assign w817[28] = |(datain[199:196] ^ 5);
  assign w817[29] = |(datain[195:192] ^ 11);
  assign w817[30] = |(datain[191:188] ^ 12);
  assign w817[31] = |(datain[187:184] ^ 3);
  assign w817[32] = |(datain[183:180] ^ 14);
  assign w817[33] = |(datain[179:176] ^ 8);
  assign w817[34] = |(datain[175:172] ^ 14);
  assign w817[35] = |(datain[171:168] ^ 2);
  assign w817[36] = |(datain[167:164] ^ 15);
  assign w817[37] = |(datain[163:160] ^ 15);
  assign w817[38] = |(datain[159:156] ^ 11);
  assign w817[39] = |(datain[155:152] ^ 4);
  assign w817[40] = |(datain[151:148] ^ 4);
  assign w817[41] = |(datain[147:144] ^ 0);
  assign w817[42] = |(datain[143:140] ^ 11);
  assign w817[43] = |(datain[139:136] ^ 9);
  assign w817[44] = |(datain[135:132] ^ 9);
  assign w817[45] = |(datain[131:128] ^ 12);
  assign w817[46] = |(datain[127:124] ^ 0);
  assign w817[47] = |(datain[123:120] ^ 13);
  assign w817[48] = |(datain[119:116] ^ 11);
  assign w817[49] = |(datain[115:112] ^ 10);
  assign w817[50] = |(datain[111:108] ^ 0);
  assign w817[51] = |(datain[107:104] ^ 3);
  assign w817[52] = |(datain[103:100] ^ 0);
  assign w817[53] = |(datain[99:96] ^ 1);
  assign w817[54] = |(datain[95:92] ^ 2);
  assign w817[55] = |(datain[91:88] ^ 11);
  assign w817[56] = |(datain[87:84] ^ 12);
  assign w817[57] = |(datain[83:80] ^ 10);
  assign w817[58] = |(datain[79:76] ^ 8);
  assign w817[59] = |(datain[75:72] ^ 11);
  assign w817[60] = |(datain[71:68] ^ 1);
  assign w817[61] = |(datain[67:64] ^ 14);
  assign w817[62] = |(datain[63:60] ^ 11);
  assign w817[63] = |(datain[59:56] ^ 4);
  assign w817[64] = |(datain[55:52] ^ 0);
  assign w817[65] = |(datain[51:48] ^ 13);
  assign w817[66] = |(datain[47:44] ^ 14);
  assign w817[67] = |(datain[43:40] ^ 8);
  assign w817[68] = |(datain[39:36] ^ 11);
  assign w817[69] = |(datain[35:32] ^ 1);
  assign w817[70] = |(datain[31:28] ^ 0);
  assign w817[71] = |(datain[27:24] ^ 1);
  assign comp[817] = ~(|w817);
  wire [44-1:0] w818;
  assign w818[0] = |(datain[311:308] ^ 8);
  assign w818[1] = |(datain[307:304] ^ 0);
  assign w818[2] = |(datain[303:300] ^ 15);
  assign w818[3] = |(datain[299:296] ^ 12);
  assign w818[4] = |(datain[295:292] ^ 3);
  assign w818[5] = |(datain[291:288] ^ 11);
  assign w818[6] = |(datain[287:284] ^ 7);
  assign w818[7] = |(datain[283:280] ^ 5);
  assign w818[8] = |(datain[279:276] ^ 0);
  assign w818[9] = |(datain[275:272] ^ 3);
  assign w818[10] = |(datain[271:268] ^ 14);
  assign w818[11] = |(datain[267:264] ^ 9);
  assign w818[12] = |(datain[263:260] ^ 1);
  assign w818[13] = |(datain[259:256] ^ 14);
  assign w818[14] = |(datain[255:252] ^ 15);
  assign w818[15] = |(datain[251:248] ^ 15);
  assign w818[16] = |(datain[247:244] ^ 3);
  assign w818[17] = |(datain[243:240] ^ 13);
  assign w818[18] = |(datain[239:236] ^ 0);
  assign w818[19] = |(datain[235:232] ^ 0);
  assign w818[20] = |(datain[231:228] ^ 3);
  assign w818[21] = |(datain[227:224] ^ 13);
  assign w818[22] = |(datain[223:220] ^ 7);
  assign w818[23] = |(datain[219:216] ^ 4);
  assign w818[24] = |(datain[215:212] ^ 0);
  assign w818[25] = |(datain[211:208] ^ 15);
  assign w818[26] = |(datain[207:204] ^ 3);
  assign w818[27] = |(datain[203:200] ^ 13);
  assign w818[28] = |(datain[199:196] ^ 0);
  assign w818[29] = |(datain[195:192] ^ 2);
  assign w818[30] = |(datain[191:188] ^ 3);
  assign w818[31] = |(datain[187:184] ^ 13);
  assign w818[32] = |(datain[183:180] ^ 7);
  assign w818[33] = |(datain[179:176] ^ 4);
  assign w818[34] = |(datain[175:172] ^ 0);
  assign w818[35] = |(datain[171:168] ^ 10);
  assign w818[36] = |(datain[167:164] ^ 8);
  assign w818[37] = |(datain[163:160] ^ 0);
  assign w818[38] = |(datain[159:156] ^ 15);
  assign w818[39] = |(datain[155:152] ^ 12);
  assign w818[40] = |(datain[151:148] ^ 5);
  assign w818[41] = |(datain[147:144] ^ 6);
  assign w818[42] = |(datain[143:140] ^ 7);
  assign w818[43] = |(datain[139:136] ^ 4);
  assign comp[818] = ~(|w818);
  wire [40-1:0] w819;
  assign w819[0] = |(datain[311:308] ^ 3);
  assign w819[1] = |(datain[307:304] ^ 11);
  assign w819[2] = |(datain[303:300] ^ 7);
  assign w819[3] = |(datain[299:296] ^ 5);
  assign w819[4] = |(datain[295:292] ^ 0);
  assign w819[5] = |(datain[291:288] ^ 3);
  assign w819[6] = |(datain[287:284] ^ 14);
  assign w819[7] = |(datain[283:280] ^ 9);
  assign w819[8] = |(datain[279:276] ^ 1);
  assign w819[9] = |(datain[275:272] ^ 7);
  assign w819[10] = |(datain[271:268] ^ 15);
  assign w819[11] = |(datain[267:264] ^ 15);
  assign w819[12] = |(datain[263:260] ^ 3);
  assign w819[13] = |(datain[259:256] ^ 13);
  assign w819[14] = |(datain[255:252] ^ 0);
  assign w819[15] = |(datain[251:248] ^ 0);
  assign w819[16] = |(datain[247:244] ^ 3);
  assign w819[17] = |(datain[243:240] ^ 13);
  assign w819[18] = |(datain[239:236] ^ 7);
  assign w819[19] = |(datain[235:232] ^ 4);
  assign w819[20] = |(datain[231:228] ^ 0);
  assign w819[21] = |(datain[227:224] ^ 15);
  assign w819[22] = |(datain[223:220] ^ 3);
  assign w819[23] = |(datain[219:216] ^ 13);
  assign w819[24] = |(datain[215:212] ^ 0);
  assign w819[25] = |(datain[211:208] ^ 2);
  assign w819[26] = |(datain[207:204] ^ 3);
  assign w819[27] = |(datain[203:200] ^ 13);
  assign w819[28] = |(datain[199:196] ^ 7);
  assign w819[29] = |(datain[195:192] ^ 4);
  assign w819[30] = |(datain[191:188] ^ 0);
  assign w819[31] = |(datain[187:184] ^ 10);
  assign w819[32] = |(datain[183:180] ^ 8);
  assign w819[33] = |(datain[179:176] ^ 0);
  assign w819[34] = |(datain[175:172] ^ 15);
  assign w819[35] = |(datain[171:168] ^ 12);
  assign w819[36] = |(datain[167:164] ^ 5);
  assign w819[37] = |(datain[163:160] ^ 6);
  assign w819[38] = |(datain[159:156] ^ 7);
  assign w819[39] = |(datain[155:152] ^ 4);
  assign comp[819] = ~(|w819);
  wire [74-1:0] w820;
  assign w820[0] = |(datain[311:308] ^ 11);
  assign w820[1] = |(datain[307:304] ^ 9);
  assign w820[2] = |(datain[303:300] ^ 10);
  assign w820[3] = |(datain[299:296] ^ 5);
  assign w820[4] = |(datain[295:292] ^ 0);
  assign w820[5] = |(datain[291:288] ^ 14);
  assign w820[6] = |(datain[287:284] ^ 2);
  assign w820[7] = |(datain[283:280] ^ 11);
  assign w820[8] = |(datain[279:276] ^ 12);
  assign w820[9] = |(datain[275:272] ^ 11);
  assign w820[10] = |(datain[271:268] ^ 2);
  assign w820[11] = |(datain[267:264] ^ 14);
  assign w820[12] = |(datain[263:260] ^ 10);
  assign w820[13] = |(datain[259:256] ^ 0);
  assign w820[14] = |(datain[255:252] ^ 13);
  assign w820[15] = |(datain[251:248] ^ 14);
  assign w820[16] = |(datain[247:244] ^ 0);
  assign w820[17] = |(datain[243:240] ^ 1);
  assign w820[18] = |(datain[239:236] ^ 2);
  assign w820[19] = |(datain[235:232] ^ 14);
  assign w820[20] = |(datain[231:228] ^ 3);
  assign w820[21] = |(datain[227:224] ^ 0);
  assign w820[22] = |(datain[223:220] ^ 0);
  assign w820[23] = |(datain[219:216] ^ 7);
  assign w820[24] = |(datain[215:212] ^ 4);
  assign w820[25] = |(datain[211:208] ^ 3);
  assign w820[26] = |(datain[207:204] ^ 14);
  assign w820[27] = |(datain[203:200] ^ 2);
  assign w820[28] = |(datain[199:196] ^ 15);
  assign w820[29] = |(datain[195:192] ^ 10);
  assign w820[30] = |(datain[191:188] ^ 9);
  assign w820[31] = |(datain[187:184] ^ 13);
  assign w820[32] = |(datain[183:180] ^ 5);
  assign w820[33] = |(datain[179:176] ^ 8);
  assign w820[34] = |(datain[175:172] ^ 5);
  assign w820[35] = |(datain[171:168] ^ 9);
  assign w820[36] = |(datain[167:164] ^ 5);
  assign w820[37] = |(datain[163:160] ^ 11);
  assign w820[38] = |(datain[159:156] ^ 12);
  assign w820[39] = |(datain[155:152] ^ 3);
  assign w820[40] = |(datain[151:148] ^ 14);
  assign w820[41] = |(datain[147:144] ^ 8);
  assign w820[42] = |(datain[143:140] ^ 14);
  assign w820[43] = |(datain[139:136] ^ 2);
  assign w820[44] = |(datain[135:132] ^ 15);
  assign w820[45] = |(datain[131:128] ^ 15);
  assign w820[46] = |(datain[127:124] ^ 11);
  assign w820[47] = |(datain[123:120] ^ 4);
  assign w820[48] = |(datain[119:116] ^ 4);
  assign w820[49] = |(datain[115:112] ^ 0);
  assign w820[50] = |(datain[111:108] ^ 11);
  assign w820[51] = |(datain[107:104] ^ 9);
  assign w820[52] = |(datain[103:100] ^ 10);
  assign w820[53] = |(datain[99:96] ^ 5);
  assign w820[54] = |(datain[95:92] ^ 0);
  assign w820[55] = |(datain[91:88] ^ 14);
  assign w820[56] = |(datain[87:84] ^ 11);
  assign w820[57] = |(datain[83:80] ^ 10);
  assign w820[58] = |(datain[79:76] ^ 0);
  assign w820[59] = |(datain[75:72] ^ 3);
  assign w820[60] = |(datain[71:68] ^ 0);
  assign w820[61] = |(datain[67:64] ^ 1);
  assign w820[62] = |(datain[63:60] ^ 2);
  assign w820[63] = |(datain[59:56] ^ 11);
  assign w820[64] = |(datain[55:52] ^ 12);
  assign w820[65] = |(datain[51:48] ^ 10);
  assign w820[66] = |(datain[47:44] ^ 8);
  assign w820[67] = |(datain[43:40] ^ 11);
  assign w820[68] = |(datain[39:36] ^ 1);
  assign w820[69] = |(datain[35:32] ^ 14);
  assign w820[70] = |(datain[31:28] ^ 11);
  assign w820[71] = |(datain[27:24] ^ 14);
  assign w820[72] = |(datain[23:20] ^ 0);
  assign w820[73] = |(datain[19:16] ^ 14);
  assign comp[820] = ~(|w820);
  wire [74-1:0] w821;
  assign w821[0] = |(datain[311:308] ^ 14);
  assign w821[1] = |(datain[307:304] ^ 4);
  assign w821[2] = |(datain[303:300] ^ 15);
  assign w821[3] = |(datain[299:296] ^ 14);
  assign w821[4] = |(datain[295:292] ^ 8);
  assign w821[5] = |(datain[291:288] ^ 11);
  assign w821[6] = |(datain[287:284] ^ 1);
  assign w821[7] = |(datain[283:280] ^ 14);
  assign w821[8] = |(datain[279:276] ^ 8);
  assign w821[9] = |(datain[275:272] ^ 12);
  assign w821[10] = |(datain[271:268] ^ 0);
  assign w821[11] = |(datain[267:264] ^ 3);
  assign w821[12] = |(datain[263:260] ^ 8);
  assign w821[13] = |(datain[259:256] ^ 11);
  assign w821[14] = |(datain[255:252] ^ 1);
  assign w821[15] = |(datain[251:248] ^ 6);
  assign w821[16] = |(datain[247:244] ^ 8);
  assign w821[17] = |(datain[243:240] ^ 14);
  assign w821[18] = |(datain[239:236] ^ 0);
  assign w821[19] = |(datain[235:232] ^ 3);
  assign w821[20] = |(datain[231:228] ^ 11);
  assign w821[21] = |(datain[227:224] ^ 4);
  assign w821[22] = |(datain[223:220] ^ 4);
  assign w821[23] = |(datain[219:216] ^ 2);
  assign w821[24] = |(datain[215:212] ^ 11);
  assign w821[25] = |(datain[211:208] ^ 0);
  assign w821[26] = |(datain[207:204] ^ 0);
  assign w821[27] = |(datain[203:200] ^ 0);
  assign w821[28] = |(datain[199:196] ^ 3);
  assign w821[29] = |(datain[195:192] ^ 3);
  assign w821[30] = |(datain[191:188] ^ 12);
  assign w821[31] = |(datain[187:184] ^ 9);
  assign w821[32] = |(datain[183:180] ^ 14);
  assign w821[33] = |(datain[179:176] ^ 8);
  assign w821[34] = |(datain[175:172] ^ 13);
  assign w821[35] = |(datain[171:168] ^ 3);
  assign w821[36] = |(datain[167:164] ^ 15);
  assign w821[37] = |(datain[163:160] ^ 14);
  assign w821[38] = |(datain[159:156] ^ 11);
  assign w821[39] = |(datain[155:152] ^ 4);
  assign w821[40] = |(datain[151:148] ^ 4);
  assign w821[41] = |(datain[147:144] ^ 0);
  assign w821[42] = |(datain[143:140] ^ 11);
  assign w821[43] = |(datain[139:136] ^ 9);
  assign w821[44] = |(datain[135:132] ^ 8);
  assign w821[45] = |(datain[131:128] ^ 8);
  assign w821[46] = |(datain[127:124] ^ 0);
  assign w821[47] = |(datain[123:120] ^ 3);
  assign w821[48] = |(datain[119:116] ^ 11);
  assign w821[49] = |(datain[115:112] ^ 10);
  assign w821[50] = |(datain[111:108] ^ 0);
  assign w821[51] = |(datain[107:104] ^ 3);
  assign w821[52] = |(datain[103:100] ^ 0);
  assign w821[53] = |(datain[99:96] ^ 1);
  assign w821[54] = |(datain[95:92] ^ 2);
  assign w821[55] = |(datain[91:88] ^ 11);
  assign w821[56] = |(datain[87:84] ^ 12);
  assign w821[57] = |(datain[83:80] ^ 10);
  assign w821[58] = |(datain[79:76] ^ 0);
  assign w821[59] = |(datain[75:72] ^ 1);
  assign w821[60] = |(datain[71:68] ^ 0);
  assign w821[61] = |(datain[67:64] ^ 14);
  assign w821[62] = |(datain[63:60] ^ 8);
  assign w821[63] = |(datain[59:56] ^ 14);
  assign w821[64] = |(datain[55:52] ^ 0);
  assign w821[65] = |(datain[51:48] ^ 3);
  assign w821[66] = |(datain[47:44] ^ 8);
  assign w821[67] = |(datain[43:40] ^ 11);
  assign w821[68] = |(datain[39:36] ^ 1);
  assign w821[69] = |(datain[35:32] ^ 14);
  assign w821[70] = |(datain[31:28] ^ 8);
  assign w821[71] = |(datain[27:24] ^ 12);
  assign w821[72] = |(datain[23:20] ^ 0);
  assign w821[73] = |(datain[19:16] ^ 3);
  assign comp[821] = ~(|w821);
  wire [76-1:0] w822;
  assign w822[0] = |(datain[311:308] ^ 0);
  assign w822[1] = |(datain[307:304] ^ 1);
  assign w822[2] = |(datain[303:300] ^ 7);
  assign w822[3] = |(datain[299:296] ^ 2);
  assign w822[4] = |(datain[295:292] ^ 2);
  assign w822[5] = |(datain[291:288] ^ 2);
  assign w822[6] = |(datain[287:284] ^ 11);
  assign w822[7] = |(datain[283:280] ^ 4);
  assign w822[8] = |(datain[279:276] ^ 3);
  assign w822[9] = |(datain[275:272] ^ 12);
  assign w822[10] = |(datain[271:268] ^ 2);
  assign w822[11] = |(datain[267:264] ^ 14);
  assign w822[12] = |(datain[263:260] ^ 8);
  assign w822[13] = |(datain[259:256] ^ 11);
  assign w822[14] = |(datain[255:252] ^ 1);
  assign w822[15] = |(datain[251:248] ^ 6);
  assign w822[16] = |(datain[247:244] ^ 3);
  assign w822[17] = |(datain[243:240] ^ 14);
  assign w822[18] = |(datain[239:236] ^ 0);
  assign w822[19] = |(datain[235:232] ^ 2);
  assign w822[20] = |(datain[231:228] ^ 3);
  assign w822[21] = |(datain[227:224] ^ 3);
  assign w822[22] = |(datain[223:220] ^ 12);
  assign w822[23] = |(datain[219:216] ^ 9);
  assign w822[24] = |(datain[215:212] ^ 14);
  assign w822[25] = |(datain[211:208] ^ 8);
  assign w822[26] = |(datain[207:204] ^ 3);
  assign w822[27] = |(datain[203:200] ^ 11);
  assign w822[28] = |(datain[199:196] ^ 0);
  assign w822[29] = |(datain[195:192] ^ 1);
  assign w822[30] = |(datain[191:188] ^ 7);
  assign w822[31] = |(datain[187:184] ^ 2);
  assign w822[32] = |(datain[183:180] ^ 1);
  assign w822[33] = |(datain[179:176] ^ 4);
  assign w822[34] = |(datain[175:172] ^ 8);
  assign w822[35] = |(datain[171:168] ^ 11);
  assign w822[36] = |(datain[167:164] ^ 13);
  assign w822[37] = |(datain[163:160] ^ 8);
  assign w822[38] = |(datain[159:156] ^ 5);
  assign w822[39] = |(datain[155:152] ^ 3);
  assign w822[40] = |(datain[151:148] ^ 11);
  assign w822[41] = |(datain[147:144] ^ 4);
  assign w822[42] = |(datain[143:140] ^ 4);
  assign w822[43] = |(datain[139:136] ^ 0);
  assign w822[44] = |(datain[135:132] ^ 11);
  assign w822[45] = |(datain[131:128] ^ 10);
  assign w822[46] = |(datain[127:124] ^ 3);
  assign w822[47] = |(datain[123:120] ^ 15);
  assign w822[48] = |(datain[119:116] ^ 0);
  assign w822[49] = |(datain[115:112] ^ 12);
  assign w822[50] = |(datain[111:108] ^ 11);
  assign w822[51] = |(datain[107:104] ^ 9);
  assign w822[52] = |(datain[103:100] ^ 2);
  assign w822[53] = |(datain[99:96] ^ 9);
  assign w822[54] = |(datain[95:92] ^ 0);
  assign w822[55] = |(datain[91:88] ^ 0);
  assign w822[56] = |(datain[87:84] ^ 14);
  assign w822[57] = |(datain[83:80] ^ 8);
  assign w822[58] = |(datain[79:76] ^ 2);
  assign w822[59] = |(datain[75:72] ^ 11);
  assign w822[60] = |(datain[71:68] ^ 0);
  assign w822[61] = |(datain[67:64] ^ 1);
  assign w822[62] = |(datain[63:60] ^ 5);
  assign w822[63] = |(datain[59:56] ^ 11);
  assign w822[64] = |(datain[55:52] ^ 11);
  assign w822[65] = |(datain[51:48] ^ 4);
  assign w822[66] = |(datain[47:44] ^ 3);
  assign w822[67] = |(datain[43:40] ^ 14);
  assign w822[68] = |(datain[39:36] ^ 14);
  assign w822[69] = |(datain[35:32] ^ 8);
  assign w822[70] = |(datain[31:28] ^ 2);
  assign w822[71] = |(datain[27:24] ^ 5);
  assign w822[72] = |(datain[23:20] ^ 0);
  assign w822[73] = |(datain[19:16] ^ 1);
  assign w822[74] = |(datain[15:12] ^ 12);
  assign w822[75] = |(datain[11:8] ^ 3);
  assign comp[822] = ~(|w822);
  wire [74-1:0] w823;
  assign w823[0] = |(datain[311:308] ^ 11);
  assign w823[1] = |(datain[307:304] ^ 10);
  assign w823[2] = |(datain[303:300] ^ 1);
  assign w823[3] = |(datain[299:296] ^ 0);
  assign w823[4] = |(datain[295:292] ^ 0);
  assign w823[5] = |(datain[291:288] ^ 8);
  assign w823[6] = |(datain[287:284] ^ 12);
  assign w823[7] = |(datain[283:280] ^ 13);
  assign w823[8] = |(datain[279:276] ^ 2);
  assign w823[9] = |(datain[275:272] ^ 1);
  assign w823[10] = |(datain[271:268] ^ 3);
  assign w823[11] = |(datain[267:264] ^ 9);
  assign w823[12] = |(datain[263:260] ^ 12);
  assign w823[13] = |(datain[259:256] ^ 8);
  assign w823[14] = |(datain[255:252] ^ 7);
  assign w823[15] = |(datain[251:248] ^ 4);
  assign w823[16] = |(datain[247:244] ^ 0);
  assign w823[17] = |(datain[243:240] ^ 4);
  assign w823[18] = |(datain[239:236] ^ 11);
  assign w823[19] = |(datain[235:232] ^ 0);
  assign w823[20] = |(datain[231:228] ^ 0);
  assign w823[21] = |(datain[227:224] ^ 4);
  assign w823[22] = |(datain[223:220] ^ 14);
  assign w823[23] = |(datain[219:216] ^ 11);
  assign w823[24] = |(datain[215:212] ^ 2);
  assign w823[25] = |(datain[211:208] ^ 6);
  assign w823[26] = |(datain[207:204] ^ 11);
  assign w823[27] = |(datain[203:200] ^ 8);
  assign w823[28] = |(datain[199:196] ^ 0);
  assign w823[29] = |(datain[195:192] ^ 0);
  assign w823[30] = |(datain[191:188] ^ 4);
  assign w823[31] = |(datain[187:184] ^ 2);
  assign w823[32] = |(datain[183:180] ^ 8);
  assign w823[33] = |(datain[179:176] ^ 9);
  assign w823[34] = |(datain[175:172] ^ 15);
  assign w823[35] = |(datain[171:168] ^ 10);
  assign w823[36] = |(datain[167:164] ^ 8);
  assign w823[37] = |(datain[163:160] ^ 9);
  assign w823[38] = |(datain[159:156] ^ 15);
  assign w823[39] = |(datain[155:152] ^ 1);
  assign w823[40] = |(datain[151:148] ^ 12);
  assign w823[41] = |(datain[147:144] ^ 13);
  assign w823[42] = |(datain[143:140] ^ 2);
  assign w823[43] = |(datain[139:136] ^ 1);
  assign w823[44] = |(datain[135:132] ^ 7);
  assign w823[45] = |(datain[131:128] ^ 3);
  assign w823[46] = |(datain[127:124] ^ 0);
  assign w823[47] = |(datain[123:120] ^ 4);
  assign w823[48] = |(datain[119:116] ^ 11);
  assign w823[49] = |(datain[115:112] ^ 0);
  assign w823[50] = |(datain[111:108] ^ 0);
  assign w823[51] = |(datain[107:104] ^ 6);
  assign w823[52] = |(datain[103:100] ^ 14);
  assign w823[53] = |(datain[99:96] ^ 11);
  assign w823[54] = |(datain[95:92] ^ 1);
  assign w823[55] = |(datain[91:88] ^ 7);
  assign w823[56] = |(datain[87:84] ^ 11);
  assign w823[57] = |(datain[83:80] ^ 4);
  assign w823[58] = |(datain[79:76] ^ 4);
  assign w823[59] = |(datain[75:72] ^ 0);
  assign w823[60] = |(datain[71:68] ^ 3);
  assign w823[61] = |(datain[67:64] ^ 1);
  assign w823[62] = |(datain[63:60] ^ 13);
  assign w823[63] = |(datain[59:56] ^ 2);
  assign w823[64] = |(datain[55:52] ^ 11);
  assign w823[65] = |(datain[51:48] ^ 9);
  assign w823[66] = |(datain[47:44] ^ 12);
  assign w823[67] = |(datain[43:40] ^ 0);
  assign w823[68] = |(datain[39:36] ^ 0);
  assign w823[69] = |(datain[35:32] ^ 11);
  assign w823[70] = |(datain[31:28] ^ 12);
  assign w823[71] = |(datain[27:24] ^ 13);
  assign w823[72] = |(datain[23:20] ^ 2);
  assign w823[73] = |(datain[19:16] ^ 1);
  assign comp[823] = ~(|w823);
  wire [42-1:0] w824;
  assign w824[0] = |(datain[311:308] ^ 5);
  assign w824[1] = |(datain[307:304] ^ 11);
  assign w824[2] = |(datain[303:300] ^ 11);
  assign w824[3] = |(datain[299:296] ^ 9);
  assign w824[4] = |(datain[295:292] ^ 6);
  assign w824[5] = |(datain[291:288] ^ 14);
  assign w824[6] = |(datain[287:284] ^ 0);
  assign w824[7] = |(datain[283:280] ^ 6);
  assign w824[8] = |(datain[279:276] ^ 8);
  assign w824[9] = |(datain[275:272] ^ 3);
  assign w824[10] = |(datain[271:268] ^ 14);
  assign w824[11] = |(datain[267:264] ^ 11);
  assign w824[12] = |(datain[263:260] ^ 0);
  assign w824[13] = |(datain[259:256] ^ 3);
  assign w824[14] = |(datain[255:252] ^ 11);
  assign w824[15] = |(datain[251:248] ^ 4);
  assign w824[16] = |(datain[247:244] ^ 1);
  assign w824[17] = |(datain[243:240] ^ 5);
  assign w824[18] = |(datain[239:236] ^ 8);
  assign w824[19] = |(datain[235:232] ^ 0);
  assign w824[20] = |(datain[231:228] ^ 14);
  assign w824[21] = |(datain[227:224] ^ 12);
  assign w824[22] = |(datain[223:220] ^ 10);
  assign w824[23] = |(datain[219:216] ^ 4);
  assign w824[24] = |(datain[215:212] ^ 4);
  assign w824[25] = |(datain[211:208] ^ 11);
  assign w824[26] = |(datain[207:204] ^ 2);
  assign w824[27] = |(datain[203:200] ^ 14);
  assign w824[28] = |(datain[199:196] ^ 3);
  assign w824[29] = |(datain[195:192] ^ 0);
  assign w824[30] = |(datain[191:188] ^ 2);
  assign w824[31] = |(datain[187:184] ^ 7);
  assign w824[32] = |(datain[183:180] ^ 14);
  assign w824[33] = |(datain[179:176] ^ 2);
  assign w824[34] = |(datain[175:172] ^ 15);
  assign w824[35] = |(datain[171:168] ^ 7);
  assign w824[36] = |(datain[167:164] ^ 14);
  assign w824[37] = |(datain[163:160] ^ 9);
  assign w824[38] = |(datain[159:156] ^ 9);
  assign w824[39] = |(datain[155:152] ^ 10);
  assign w824[40] = |(datain[151:148] ^ 15);
  assign w824[41] = |(datain[147:144] ^ 9);
  assign comp[824] = ~(|w824);
  wire [32-1:0] w825;
  assign w825[0] = |(datain[311:308] ^ 0);
  assign w825[1] = |(datain[307:304] ^ 3);
  assign w825[2] = |(datain[303:300] ^ 11);
  assign w825[3] = |(datain[299:296] ^ 14);
  assign w825[4] = |(datain[295:292] ^ 0);
  assign w825[5] = |(datain[291:288] ^ 3);
  assign w825[6] = |(datain[287:284] ^ 0);
  assign w825[7] = |(datain[283:280] ^ 0);
  assign w825[8] = |(datain[279:276] ^ 11);
  assign w825[9] = |(datain[275:272] ^ 8);
  assign w825[10] = |(datain[271:268] ^ 2);
  assign w825[11] = |(datain[267:264] ^ 1);
  assign w825[12] = |(datain[263:260] ^ 3);
  assign w825[13] = |(datain[259:256] ^ 5);
  assign w825[14] = |(datain[255:252] ^ 12);
  assign w825[15] = |(datain[251:248] ^ 13);
  assign w825[16] = |(datain[247:244] ^ 2);
  assign w825[17] = |(datain[243:240] ^ 1);
  assign w825[18] = |(datain[239:236] ^ 11);
  assign w825[19] = |(datain[235:232] ^ 15);
  assign w825[20] = |(datain[231:228] ^ 0);
  assign w825[21] = |(datain[227:224] ^ 12);
  assign w825[22] = |(datain[223:220] ^ 0);
  assign w825[23] = |(datain[219:216] ^ 1);
  assign w825[24] = |(datain[215:212] ^ 0);
  assign w825[25] = |(datain[211:208] ^ 3);
  assign w825[26] = |(datain[207:204] ^ 15);
  assign w825[27] = |(datain[203:200] ^ 14);
  assign w825[28] = |(datain[199:196] ^ 2);
  assign w825[29] = |(datain[195:192] ^ 14);
  assign w825[30] = |(datain[191:188] ^ 8);
  assign w825[31] = |(datain[187:184] ^ 9);
  assign comp[825] = ~(|w825);
  wire [28-1:0] w826;
  assign w826[0] = |(datain[311:308] ^ 0);
  assign w826[1] = |(datain[307:304] ^ 2);
  assign w826[2] = |(datain[303:300] ^ 7);
  assign w826[3] = |(datain[299:296] ^ 2);
  assign w826[4] = |(datain[295:292] ^ 0);
  assign w826[5] = |(datain[291:288] ^ 13);
  assign w826[6] = |(datain[287:284] ^ 8);
  assign w826[7] = |(datain[283:280] ^ 0);
  assign w826[8] = |(datain[279:276] ^ 15);
  assign w826[9] = |(datain[275:272] ^ 12);
  assign w826[10] = |(datain[271:268] ^ 0);
  assign w826[11] = |(datain[267:264] ^ 4);
  assign w826[12] = |(datain[263:260] ^ 7);
  assign w826[13] = |(datain[259:256] ^ 3);
  assign w826[14] = |(datain[255:252] ^ 0);
  assign w826[15] = |(datain[251:248] ^ 8);
  assign w826[16] = |(datain[247:244] ^ 8);
  assign w826[17] = |(datain[243:240] ^ 0);
  assign w826[18] = |(datain[239:236] ^ 15);
  assign w826[19] = |(datain[235:232] ^ 10);
  assign w826[20] = |(datain[231:228] ^ 8);
  assign w826[21] = |(datain[227:224] ^ 0);
  assign w826[22] = |(datain[223:220] ^ 7);
  assign w826[23] = |(datain[219:216] ^ 3);
  assign w826[24] = |(datain[215:212] ^ 0);
  assign w826[25] = |(datain[211:208] ^ 3);
  assign w826[26] = |(datain[207:204] ^ 14);
  assign w826[27] = |(datain[203:200] ^ 8);
  assign comp[826] = ~(|w826);
  wire [42-1:0] w827;
  assign w827[0] = |(datain[311:308] ^ 11);
  assign w827[1] = |(datain[307:304] ^ 11);
  assign w827[2] = |(datain[303:300] ^ 0);
  assign w827[3] = |(datain[299:296] ^ 2);
  assign w827[4] = |(datain[295:292] ^ 0);
  assign w827[5] = |(datain[291:288] ^ 1);
  assign w827[6] = |(datain[287:284] ^ 12);
  assign w827[7] = |(datain[283:280] ^ 13);
  assign w827[8] = |(datain[279:276] ^ 2);
  assign w827[9] = |(datain[275:272] ^ 1);
  assign w827[10] = |(datain[271:268] ^ 8);
  assign w827[11] = |(datain[267:264] ^ 6);
  assign w827[12] = |(datain[263:260] ^ 15);
  assign w827[13] = |(datain[259:256] ^ 11);
  assign w827[14] = |(datain[255:252] ^ 3);
  assign w827[15] = |(datain[251:248] ^ 11);
  assign w827[16] = |(datain[247:244] ^ 12);
  assign w827[17] = |(datain[243:240] ^ 3);
  assign w827[18] = |(datain[239:236] ^ 7);
  assign w827[19] = |(datain[235:232] ^ 5);
  assign w827[20] = |(datain[231:228] ^ 0);
  assign w827[21] = |(datain[227:224] ^ 2);
  assign w827[22] = |(datain[223:220] ^ 14);
  assign w827[23] = |(datain[219:216] ^ 11);
  assign w827[24] = |(datain[215:212] ^ 6);
  assign w827[25] = |(datain[211:208] ^ 3);
  assign w827[26] = |(datain[207:204] ^ 1);
  assign w827[27] = |(datain[203:200] ^ 14);
  assign w827[28] = |(datain[199:196] ^ 5);
  assign w827[29] = |(datain[195:192] ^ 8);
  assign w827[30] = |(datain[191:188] ^ 2);
  assign w827[31] = |(datain[187:184] ^ 13);
  assign w827[32] = |(datain[183:180] ^ 0);
  assign w827[33] = |(datain[179:176] ^ 4);
  assign w827[34] = |(datain[175:172] ^ 0);
  assign w827[35] = |(datain[171:168] ^ 0);
  assign w827[36] = |(datain[167:164] ^ 8);
  assign w827[37] = |(datain[163:160] ^ 14);
  assign w827[38] = |(datain[159:156] ^ 12);
  assign w827[39] = |(datain[155:152] ^ 0);
  assign w827[40] = |(datain[151:148] ^ 2);
  assign w827[41] = |(datain[147:144] ^ 6);
  assign comp[827] = ~(|w827);
  wire [76-1:0] w828;
  assign w828[0] = |(datain[311:308] ^ 13);
  assign w828[1] = |(datain[307:304] ^ 12);
  assign w828[2] = |(datain[303:300] ^ 0);
  assign w828[3] = |(datain[299:296] ^ 0);
  assign w828[4] = |(datain[295:292] ^ 1);
  assign w828[5] = |(datain[291:288] ^ 13);
  assign w828[6] = |(datain[287:284] ^ 10);
  assign w828[7] = |(datain[283:280] ^ 12);
  assign w828[8] = |(datain[279:276] ^ 14);
  assign w828[9] = |(datain[275:272] ^ 8);
  assign w828[10] = |(datain[271:268] ^ 8);
  assign w828[11] = |(datain[267:264] ^ 1);
  assign w828[12] = |(datain[263:260] ^ 15);
  assign w828[13] = |(datain[259:256] ^ 14);
  assign w828[14] = |(datain[255:252] ^ 11);
  assign w828[15] = |(datain[251:248] ^ 4);
  assign w828[16] = |(datain[247:244] ^ 4);
  assign w828[17] = |(datain[243:240] ^ 0);
  assign w828[18] = |(datain[239:236] ^ 11);
  assign w828[19] = |(datain[235:232] ^ 9);
  assign w828[20] = |(datain[231:228] ^ 6);
  assign w828[21] = |(datain[227:224] ^ 5);
  assign w828[22] = |(datain[223:220] ^ 0);
  assign w828[23] = |(datain[219:216] ^ 3);
  assign w828[24] = |(datain[215:212] ^ 0);
  assign w828[25] = |(datain[211:208] ^ 14);
  assign w828[26] = |(datain[207:204] ^ 1);
  assign w828[27] = |(datain[203:200] ^ 15);
  assign w828[28] = |(datain[199:196] ^ 11);
  assign w828[29] = |(datain[195:192] ^ 10);
  assign w828[30] = |(datain[191:188] ^ 6);
  assign w828[31] = |(datain[187:184] ^ 7);
  assign w828[32] = |(datain[183:180] ^ 0);
  assign w828[33] = |(datain[179:176] ^ 3);
  assign w828[34] = |(datain[175:172] ^ 12);
  assign w828[35] = |(datain[171:168] ^ 12);
  assign w828[36] = |(datain[167:164] ^ 7);
  assign w828[37] = |(datain[163:160] ^ 2);
  assign w828[38] = |(datain[159:156] ^ 2);
  assign w828[39] = |(datain[155:152] ^ 1);
  assign w828[40] = |(datain[151:148] ^ 11);
  assign w828[41] = |(datain[147:144] ^ 8);
  assign w828[42] = |(datain[143:140] ^ 0);
  assign w828[43] = |(datain[139:136] ^ 0);
  assign w828[44] = |(datain[135:132] ^ 4);
  assign w828[45] = |(datain[131:128] ^ 2);
  assign w828[46] = |(datain[127:124] ^ 3);
  assign w828[47] = |(datain[123:120] ^ 3);
  assign w828[48] = |(datain[119:116] ^ 12);
  assign w828[49] = |(datain[115:112] ^ 9);
  assign w828[50] = |(datain[111:108] ^ 3);
  assign w828[51] = |(datain[107:104] ^ 3);
  assign w828[52] = |(datain[103:100] ^ 13);
  assign w828[53] = |(datain[99:96] ^ 2);
  assign w828[54] = |(datain[95:92] ^ 12);
  assign w828[55] = |(datain[91:88] ^ 12);
  assign w828[56] = |(datain[87:84] ^ 11);
  assign w828[57] = |(datain[83:80] ^ 4);
  assign w828[58] = |(datain[79:76] ^ 4);
  assign w828[59] = |(datain[75:72] ^ 0);
  assign w828[60] = |(datain[71:68] ^ 11);
  assign w828[61] = |(datain[67:64] ^ 9);
  assign w828[62] = |(datain[63:60] ^ 1);
  assign w828[63] = |(datain[59:56] ^ 8);
  assign w828[64] = |(datain[55:52] ^ 0);
  assign w828[65] = |(datain[51:48] ^ 0);
  assign w828[66] = |(datain[47:44] ^ 11);
  assign w828[67] = |(datain[43:40] ^ 10);
  assign w828[68] = |(datain[39:36] ^ 12);
  assign w828[69] = |(datain[35:32] ^ 10);
  assign w828[70] = |(datain[31:28] ^ 0);
  assign w828[71] = |(datain[27:24] ^ 0);
  assign w828[72] = |(datain[23:20] ^ 12);
  assign w828[73] = |(datain[19:16] ^ 12);
  assign w828[74] = |(datain[15:12] ^ 7);
  assign w828[75] = |(datain[11:8] ^ 2);
  assign comp[828] = ~(|w828);
  wire [74-1:0] w829;
  assign w829[0] = |(datain[311:308] ^ 10);
  assign w829[1] = |(datain[307:304] ^ 3);
  assign w829[2] = |(datain[303:300] ^ 9);
  assign w829[3] = |(datain[299:296] ^ 15);
  assign w829[4] = |(datain[295:292] ^ 0);
  assign w829[5] = |(datain[291:288] ^ 1);
  assign w829[6] = |(datain[287:284] ^ 11);
  assign w829[7] = |(datain[283:280] ^ 10);
  assign w829[8] = |(datain[279:276] ^ 11);
  assign w829[9] = |(datain[275:272] ^ 2);
  assign w829[10] = |(datain[271:268] ^ 0);
  assign w829[11] = |(datain[267:264] ^ 3);
  assign w829[12] = |(datain[263:260] ^ 11);
  assign w829[13] = |(datain[259:256] ^ 9);
  assign w829[14] = |(datain[255:252] ^ 11);
  assign w829[15] = |(datain[251:248] ^ 2);
  assign w829[16] = |(datain[247:244] ^ 0);
  assign w829[17] = |(datain[243:240] ^ 1);
  assign w829[18] = |(datain[239:236] ^ 11);
  assign w829[19] = |(datain[235:232] ^ 4);
  assign w829[20] = |(datain[231:228] ^ 4);
  assign w829[21] = |(datain[227:224] ^ 0);
  assign w829[22] = |(datain[223:220] ^ 12);
  assign w829[23] = |(datain[219:216] ^ 13);
  assign w829[24] = |(datain[215:212] ^ 2);
  assign w829[25] = |(datain[211:208] ^ 1);
  assign w829[26] = |(datain[207:204] ^ 12);
  assign w829[27] = |(datain[203:200] ^ 6);
  assign w829[28] = |(datain[199:196] ^ 0);
  assign w829[29] = |(datain[195:192] ^ 6);
  assign w829[30] = |(datain[191:188] ^ 1);
  assign w829[31] = |(datain[187:184] ^ 2);
  assign w829[32] = |(datain[183:180] ^ 0);
  assign w829[33] = |(datain[179:176] ^ 2);
  assign w829[34] = |(datain[175:172] ^ 4);
  assign w829[35] = |(datain[171:168] ^ 14);
  assign w829[36] = |(datain[167:164] ^ 11);
  assign w829[37] = |(datain[163:160] ^ 8);
  assign w829[38] = |(datain[159:156] ^ 0);
  assign w829[39] = |(datain[155:152] ^ 0);
  assign w829[40] = |(datain[151:148] ^ 4);
  assign w829[41] = |(datain[147:144] ^ 2);
  assign w829[42] = |(datain[143:140] ^ 3);
  assign w829[43] = |(datain[139:136] ^ 3);
  assign w829[44] = |(datain[135:132] ^ 12);
  assign w829[45] = |(datain[131:128] ^ 9);
  assign w829[46] = |(datain[127:124] ^ 3);
  assign w829[47] = |(datain[123:120] ^ 3);
  assign w829[48] = |(datain[119:116] ^ 13);
  assign w829[49] = |(datain[115:112] ^ 2);
  assign w829[50] = |(datain[111:108] ^ 12);
  assign w829[51] = |(datain[107:104] ^ 13);
  assign w829[52] = |(datain[103:100] ^ 2);
  assign w829[53] = |(datain[99:96] ^ 1);
  assign w829[54] = |(datain[95:92] ^ 11);
  assign w829[55] = |(datain[91:88] ^ 4);
  assign w829[56] = |(datain[87:84] ^ 4);
  assign w829[57] = |(datain[83:80] ^ 0);
  assign w829[58] = |(datain[79:76] ^ 11);
  assign w829[59] = |(datain[75:72] ^ 10);
  assign w829[60] = |(datain[71:68] ^ 0);
  assign w829[61] = |(datain[67:64] ^ 0);
  assign w829[62] = |(datain[63:60] ^ 0);
  assign w829[63] = |(datain[59:56] ^ 1);
  assign w829[64] = |(datain[55:52] ^ 11);
  assign w829[65] = |(datain[51:48] ^ 9);
  assign w829[66] = |(datain[47:44] ^ 11);
  assign w829[67] = |(datain[43:40] ^ 2);
  assign w829[68] = |(datain[39:36] ^ 0);
  assign w829[69] = |(datain[35:32] ^ 1);
  assign w829[70] = |(datain[31:28] ^ 12);
  assign w829[71] = |(datain[27:24] ^ 13);
  assign w829[72] = |(datain[23:20] ^ 2);
  assign w829[73] = |(datain[19:16] ^ 1);
  assign comp[829] = ~(|w829);
  wire [74-1:0] w830;
  assign w830[0] = |(datain[311:308] ^ 11);
  assign w830[1] = |(datain[307:304] ^ 10);
  assign w830[2] = |(datain[303:300] ^ 6);
  assign w830[3] = |(datain[299:296] ^ 8);
  assign w830[4] = |(datain[295:292] ^ 0);
  assign w830[5] = |(datain[291:288] ^ 1);
  assign w830[6] = |(datain[287:284] ^ 11);
  assign w830[7] = |(datain[283:280] ^ 4);
  assign w830[8] = |(datain[279:276] ^ 4);
  assign w830[9] = |(datain[275:272] ^ 0);
  assign w830[10] = |(datain[271:268] ^ 12);
  assign w830[11] = |(datain[267:264] ^ 13);
  assign w830[12] = |(datain[263:260] ^ 2);
  assign w830[13] = |(datain[259:256] ^ 1);
  assign w830[14] = |(datain[255:252] ^ 11);
  assign w830[15] = |(datain[251:248] ^ 0);
  assign w830[16] = |(datain[247:244] ^ 0);
  assign w830[17] = |(datain[243:240] ^ 2);
  assign w830[18] = |(datain[239:236] ^ 3);
  assign w830[19] = |(datain[235:232] ^ 3);
  assign w830[20] = |(datain[231:228] ^ 13);
  assign w830[21] = |(datain[227:224] ^ 2);
  assign w830[22] = |(datain[223:220] ^ 3);
  assign w830[23] = |(datain[219:216] ^ 3);
  assign w830[24] = |(datain[215:212] ^ 12);
  assign w830[25] = |(datain[211:208] ^ 9);
  assign w830[26] = |(datain[207:204] ^ 14);
  assign w830[27] = |(datain[203:200] ^ 8);
  assign w830[28] = |(datain[199:196] ^ 7);
  assign w830[29] = |(datain[195:192] ^ 7);
  assign w830[30] = |(datain[191:188] ^ 0);
  assign w830[31] = |(datain[187:184] ^ 0);
  assign w830[32] = |(datain[183:180] ^ 11);
  assign w830[33] = |(datain[179:176] ^ 4);
  assign w830[34] = |(datain[175:172] ^ 4);
  assign w830[35] = |(datain[171:168] ^ 0);
  assign w830[36] = |(datain[167:164] ^ 11);
  assign w830[37] = |(datain[163:160] ^ 9);
  assign w830[38] = |(datain[159:156] ^ 4);
  assign w830[39] = |(datain[155:152] ^ 9);
  assign w830[40] = |(datain[151:148] ^ 0);
  assign w830[41] = |(datain[147:144] ^ 2);
  assign w830[42] = |(datain[143:140] ^ 11);
  assign w830[43] = |(datain[139:136] ^ 10);
  assign w830[44] = |(datain[135:132] ^ 0);
  assign w830[45] = |(datain[131:128] ^ 0);
  assign w830[46] = |(datain[127:124] ^ 0);
  assign w830[47] = |(datain[123:120] ^ 1);
  assign w830[48] = |(datain[119:116] ^ 12);
  assign w830[49] = |(datain[115:112] ^ 13);
  assign w830[50] = |(datain[111:108] ^ 2);
  assign w830[51] = |(datain[107:104] ^ 1);
  assign w830[52] = |(datain[103:100] ^ 11);
  assign w830[53] = |(datain[99:96] ^ 8);
  assign w830[54] = |(datain[95:92] ^ 0);
  assign w830[55] = |(datain[91:88] ^ 0);
  assign w830[56] = |(datain[87:84] ^ 3);
  assign w830[57] = |(datain[83:80] ^ 14);
  assign w830[58] = |(datain[79:76] ^ 12);
  assign w830[59] = |(datain[75:72] ^ 13);
  assign w830[60] = |(datain[71:68] ^ 2);
  assign w830[61] = |(datain[67:64] ^ 1);
  assign w830[62] = |(datain[63:60] ^ 1);
  assign w830[63] = |(datain[59:56] ^ 15);
  assign w830[64] = |(datain[55:52] ^ 5);
  assign w830[65] = |(datain[51:48] ^ 10);
  assign w830[66] = |(datain[47:44] ^ 5);
  assign w830[67] = |(datain[43:40] ^ 9);
  assign w830[68] = |(datain[39:36] ^ 14);
  assign w830[69] = |(datain[35:32] ^ 8);
  assign w830[70] = |(datain[31:28] ^ 12);
  assign w830[71] = |(datain[27:24] ^ 0);
  assign w830[72] = |(datain[23:20] ^ 0);
  assign w830[73] = |(datain[19:16] ^ 0);
  assign comp[830] = ~(|w830);
  wire [76-1:0] w831;
  assign w831[0] = |(datain[311:308] ^ 11);
  assign w831[1] = |(datain[307:304] ^ 0);
  assign w831[2] = |(datain[303:300] ^ 4);
  assign w831[3] = |(datain[299:296] ^ 0);
  assign w831[4] = |(datain[295:292] ^ 3);
  assign w831[5] = |(datain[291:288] ^ 3);
  assign w831[6] = |(datain[287:284] ^ 12);
  assign w831[7] = |(datain[283:280] ^ 9);
  assign w831[8] = |(datain[279:276] ^ 0);
  assign w831[9] = |(datain[275:272] ^ 5);
  assign w831[10] = |(datain[271:268] ^ 0);
  assign w831[11] = |(datain[267:264] ^ 0);
  assign w831[12] = |(datain[263:260] ^ 0);
  assign w831[13] = |(datain[259:256] ^ 1);
  assign w831[14] = |(datain[255:252] ^ 4);
  assign w831[15] = |(datain[251:248] ^ 0);
  assign w831[16] = |(datain[247:244] ^ 0);
  assign w831[17] = |(datain[243:240] ^ 5);
  assign w831[18] = |(datain[239:236] ^ 4);
  assign w831[19] = |(datain[235:232] ^ 14);
  assign w831[20] = |(datain[231:228] ^ 0);
  assign w831[21] = |(datain[227:224] ^ 0);
  assign w831[22] = |(datain[223:220] ^ 4);
  assign w831[23] = |(datain[219:216] ^ 0);
  assign w831[24] = |(datain[215:212] ^ 12);
  assign w831[25] = |(datain[211:208] ^ 13);
  assign w831[26] = |(datain[207:204] ^ 2);
  assign w831[27] = |(datain[203:200] ^ 1);
  assign w831[28] = |(datain[199:196] ^ 5);
  assign w831[29] = |(datain[195:192] ^ 0);
  assign w831[30] = |(datain[191:188] ^ 1);
  assign w831[31] = |(datain[187:184] ^ 14);
  assign w831[32] = |(datain[183:180] ^ 5);
  assign w831[33] = |(datain[179:176] ^ 1);
  assign w831[34] = |(datain[175:172] ^ 5);
  assign w831[35] = |(datain[171:168] ^ 9);
  assign w831[36] = |(datain[167:164] ^ 1);
  assign w831[37] = |(datain[163:160] ^ 15);
  assign w831[38] = |(datain[159:156] ^ 5);
  assign w831[39] = |(datain[155:152] ^ 8);
  assign w831[40] = |(datain[151:148] ^ 11);
  assign w831[41] = |(datain[147:144] ^ 4);
  assign w831[42] = |(datain[143:140] ^ 2);
  assign w831[43] = |(datain[139:136] ^ 0);
  assign w831[44] = |(datain[135:132] ^ 8);
  assign w831[45] = |(datain[131:128] ^ 0);
  assign w831[46] = |(datain[127:124] ^ 12);
  assign w831[47] = |(datain[123:120] ^ 4);
  assign w831[48] = |(datain[119:116] ^ 1);
  assign w831[49] = |(datain[115:112] ^ 5);
  assign w831[50] = |(datain[111:108] ^ 8);
  assign w831[51] = |(datain[107:104] ^ 0);
  assign w831[52] = |(datain[103:100] ^ 12);
  assign w831[53] = |(datain[99:96] ^ 4);
  assign w831[54] = |(datain[95:92] ^ 0);
  assign w831[55] = |(datain[91:88] ^ 10);
  assign w831[56] = |(datain[87:84] ^ 15);
  assign w831[57] = |(datain[83:80] ^ 14);
  assign w831[58] = |(datain[79:76] ^ 12);
  assign w831[59] = |(datain[75:72] ^ 4);
  assign w831[60] = |(datain[71:68] ^ 11);
  assign w831[61] = |(datain[67:64] ^ 9);
  assign w831[62] = |(datain[63:60] ^ 1);
  assign w831[63] = |(datain[59:56] ^ 10);
  assign w831[64] = |(datain[55:52] ^ 0);
  assign w831[65] = |(datain[51:48] ^ 0);
  assign w831[66] = |(datain[47:44] ^ 11);
  assign w831[67] = |(datain[43:40] ^ 10);
  assign w831[68] = |(datain[39:36] ^ 11);
  assign w831[69] = |(datain[35:32] ^ 1);
  assign w831[70] = |(datain[31:28] ^ 0);
  assign w831[71] = |(datain[27:24] ^ 2);
  assign w831[72] = |(datain[23:20] ^ 12);
  assign w831[73] = |(datain[19:16] ^ 13);
  assign w831[74] = |(datain[15:12] ^ 2);
  assign w831[75] = |(datain[11:8] ^ 1);
  assign comp[831] = ~(|w831);
  wire [74-1:0] w832;
  assign w832[0] = |(datain[311:308] ^ 3);
  assign w832[1] = |(datain[307:304] ^ 3);
  assign w832[2] = |(datain[303:300] ^ 12);
  assign w832[3] = |(datain[299:296] ^ 9);
  assign w832[4] = |(datain[295:292] ^ 0);
  assign w832[5] = |(datain[291:288] ^ 5);
  assign w832[6] = |(datain[287:284] ^ 0);
  assign w832[7] = |(datain[283:280] ^ 0);
  assign w832[8] = |(datain[279:276] ^ 0);
  assign w832[9] = |(datain[275:272] ^ 1);
  assign w832[10] = |(datain[271:268] ^ 4);
  assign w832[11] = |(datain[267:264] ^ 0);
  assign w832[12] = |(datain[263:260] ^ 0);
  assign w832[13] = |(datain[259:256] ^ 5);
  assign w832[14] = |(datain[255:252] ^ 4);
  assign w832[15] = |(datain[251:248] ^ 14);
  assign w832[16] = |(datain[247:244] ^ 0);
  assign w832[17] = |(datain[243:240] ^ 0);
  assign w832[18] = |(datain[239:236] ^ 4);
  assign w832[19] = |(datain[235:232] ^ 0);
  assign w832[20] = |(datain[231:228] ^ 12);
  assign w832[21] = |(datain[227:224] ^ 13);
  assign w832[22] = |(datain[223:220] ^ 2);
  assign w832[23] = |(datain[219:216] ^ 1);
  assign w832[24] = |(datain[215:212] ^ 5);
  assign w832[25] = |(datain[211:208] ^ 0);
  assign w832[26] = |(datain[207:204] ^ 1);
  assign w832[27] = |(datain[203:200] ^ 14);
  assign w832[28] = |(datain[199:196] ^ 5);
  assign w832[29] = |(datain[195:192] ^ 1);
  assign w832[30] = |(datain[191:188] ^ 5);
  assign w832[31] = |(datain[187:184] ^ 9);
  assign w832[32] = |(datain[183:180] ^ 1);
  assign w832[33] = |(datain[179:176] ^ 15);
  assign w832[34] = |(datain[175:172] ^ 5);
  assign w832[35] = |(datain[171:168] ^ 8);
  assign w832[36] = |(datain[167:164] ^ 11);
  assign w832[37] = |(datain[163:160] ^ 4);
  assign w832[38] = |(datain[159:156] ^ 2);
  assign w832[39] = |(datain[155:152] ^ 0);
  assign w832[40] = |(datain[151:148] ^ 8);
  assign w832[41] = |(datain[147:144] ^ 0);
  assign w832[42] = |(datain[143:140] ^ 12);
  assign w832[43] = |(datain[139:136] ^ 4);
  assign w832[44] = |(datain[135:132] ^ 1);
  assign w832[45] = |(datain[131:128] ^ 5);
  assign w832[46] = |(datain[127:124] ^ 8);
  assign w832[47] = |(datain[123:120] ^ 0);
  assign w832[48] = |(datain[119:116] ^ 12);
  assign w832[49] = |(datain[115:112] ^ 4);
  assign w832[50] = |(datain[111:108] ^ 0);
  assign w832[51] = |(datain[107:104] ^ 10);
  assign w832[52] = |(datain[103:100] ^ 15);
  assign w832[53] = |(datain[99:96] ^ 14);
  assign w832[54] = |(datain[95:92] ^ 12);
  assign w832[55] = |(datain[91:88] ^ 4);
  assign w832[56] = |(datain[87:84] ^ 11);
  assign w832[57] = |(datain[83:80] ^ 9);
  assign w832[58] = |(datain[79:76] ^ 1);
  assign w832[59] = |(datain[75:72] ^ 10);
  assign w832[60] = |(datain[71:68] ^ 0);
  assign w832[61] = |(datain[67:64] ^ 0);
  assign w832[62] = |(datain[63:60] ^ 11);
  assign w832[63] = |(datain[59:56] ^ 10);
  assign w832[64] = |(datain[55:52] ^ 10);
  assign w832[65] = |(datain[51:48] ^ 10);
  assign w832[66] = |(datain[47:44] ^ 0);
  assign w832[67] = |(datain[43:40] ^ 2);
  assign w832[68] = |(datain[39:36] ^ 12);
  assign w832[69] = |(datain[35:32] ^ 13);
  assign w832[70] = |(datain[31:28] ^ 2);
  assign w832[71] = |(datain[27:24] ^ 1);
  assign w832[72] = |(datain[23:20] ^ 5);
  assign w832[73] = |(datain[19:16] ^ 2);
  assign comp[832] = ~(|w832);
  wire [32-1:0] w833;
  assign w833[0] = |(datain[311:308] ^ 11);
  assign w833[1] = |(datain[307:304] ^ 4);
  assign w833[2] = |(datain[303:300] ^ 15);
  assign w833[3] = |(datain[299:296] ^ 15);
  assign w833[4] = |(datain[295:292] ^ 12);
  assign w833[5] = |(datain[291:288] ^ 13);
  assign w833[6] = |(datain[287:284] ^ 2);
  assign w833[7] = |(datain[283:280] ^ 1);
  assign w833[8] = |(datain[279:276] ^ 8);
  assign w833[9] = |(datain[275:272] ^ 0);
  assign w833[10] = |(datain[271:268] ^ 15);
  assign w833[11] = |(datain[267:264] ^ 12);
  assign w833[12] = |(datain[263:260] ^ 15);
  assign w833[13] = |(datain[259:256] ^ 10);
  assign w833[14] = |(datain[255:252] ^ 7);
  assign w833[15] = |(datain[251:248] ^ 5);
  assign w833[16] = |(datain[247:244] ^ 0);
  assign w833[17] = |(datain[243:240] ^ 3);
  assign w833[18] = |(datain[239:236] ^ 14);
  assign w833[19] = |(datain[235:232] ^ 11);
  assign w833[20] = |(datain[231:228] ^ 6);
  assign w833[21] = |(datain[227:224] ^ 1);
  assign w833[22] = |(datain[223:220] ^ 9);
  assign w833[23] = |(datain[219:216] ^ 0);
  assign w833[24] = |(datain[215:212] ^ 1);
  assign w833[25] = |(datain[211:208] ^ 14);
  assign w833[26] = |(datain[207:204] ^ 3);
  assign w833[27] = |(datain[203:200] ^ 1);
  assign w833[28] = |(datain[199:196] ^ 12);
  assign w833[29] = |(datain[195:192] ^ 0);
  assign w833[30] = |(datain[191:188] ^ 8);
  assign w833[31] = |(datain[187:184] ^ 14);
  assign comp[833] = ~(|w833);
  wire [42-1:0] w834;
  assign w834[0] = |(datain[311:308] ^ 3);
  assign w834[1] = |(datain[307:304] ^ 1);
  assign w834[2] = |(datain[303:300] ^ 12);
  assign w834[3] = |(datain[299:296] ^ 9);
  assign w834[4] = |(datain[295:292] ^ 3);
  assign w834[5] = |(datain[291:288] ^ 1);
  assign w834[6] = |(datain[287:284] ^ 13);
  assign w834[7] = |(datain[283:280] ^ 2);
  assign w834[8] = |(datain[279:276] ^ 14);
  assign w834[9] = |(datain[275:272] ^ 8);
  assign w834[10] = |(datain[271:268] ^ 4);
  assign w834[11] = |(datain[267:264] ^ 5);
  assign w834[12] = |(datain[263:260] ^ 0);
  assign w834[13] = |(datain[259:256] ^ 0);
  assign w834[14] = |(datain[255:252] ^ 11);
  assign w834[15] = |(datain[251:248] ^ 4);
  assign w834[16] = |(datain[247:244] ^ 4);
  assign w834[17] = |(datain[243:240] ^ 0);
  assign w834[18] = |(datain[239:236] ^ 12);
  assign w834[19] = |(datain[235:232] ^ 7);
  assign w834[20] = |(datain[231:228] ^ 12);
  assign w834[21] = |(datain[227:224] ^ 2);
  assign w834[22] = |(datain[223:220] ^ 0);
  assign w834[23] = |(datain[219:216] ^ 0);
  assign w834[24] = |(datain[215:212] ^ 0);
  assign w834[25] = |(datain[211:208] ^ 5);
  assign w834[26] = |(datain[207:204] ^ 5);
  assign w834[27] = |(datain[203:200] ^ 9);
  assign w834[28] = |(datain[199:196] ^ 8);
  assign w834[29] = |(datain[195:192] ^ 1);
  assign w834[30] = |(datain[191:188] ^ 12);
  assign w834[31] = |(datain[187:184] ^ 1);
  assign w834[32] = |(datain[183:180] ^ 0);
  assign w834[33] = |(datain[179:176] ^ 0);
  assign w834[34] = |(datain[175:172] ^ 0);
  assign w834[35] = |(datain[171:168] ^ 4);
  assign w834[36] = |(datain[167:164] ^ 14);
  assign w834[37] = |(datain[163:160] ^ 8);
  assign w834[38] = |(datain[159:156] ^ 3);
  assign w834[39] = |(datain[155:152] ^ 7);
  assign w834[40] = |(datain[151:148] ^ 0);
  assign w834[41] = |(datain[147:144] ^ 0);
  assign comp[834] = ~(|w834);
  wire [50-1:0] w835;
  assign w835[0] = |(datain[311:308] ^ 0);
  assign w835[1] = |(datain[307:304] ^ 3);
  assign w835[2] = |(datain[303:300] ^ 0);
  assign w835[3] = |(datain[299:296] ^ 1);
  assign w835[4] = |(datain[295:292] ^ 8);
  assign w835[5] = |(datain[291:288] ^ 13);
  assign w835[6] = |(datain[287:284] ^ 9);
  assign w835[7] = |(datain[283:280] ^ 14);
  assign w835[8] = |(datain[279:276] ^ 2);
  assign w835[9] = |(datain[275:272] ^ 0);
  assign w835[10] = |(datain[271:268] ^ 0);
  assign w835[11] = |(datain[267:264] ^ 1);
  assign w835[12] = |(datain[263:260] ^ 8);
  assign w835[13] = |(datain[259:256] ^ 13);
  assign w835[14] = |(datain[255:252] ^ 9);
  assign w835[15] = |(datain[251:248] ^ 6);
  assign w835[16] = |(datain[247:244] ^ 8);
  assign w835[17] = |(datain[243:240] ^ 11);
  assign w835[18] = |(datain[239:236] ^ 0);
  assign w835[19] = |(datain[235:232] ^ 1);
  assign w835[20] = |(datain[231:228] ^ 3);
  assign w835[21] = |(datain[227:224] ^ 14);
  assign w835[22] = |(datain[223:220] ^ 8);
  assign w835[23] = |(datain[219:216] ^ 10);
  assign w835[24] = |(datain[215:212] ^ 8);
  assign w835[25] = |(datain[211:208] ^ 14);
  assign w835[26] = |(datain[207:204] ^ 0);
  assign w835[27] = |(datain[203:200] ^ 3);
  assign w835[28] = |(datain[199:196] ^ 0);
  assign w835[29] = |(datain[195:192] ^ 1);
  assign w835[30] = |(datain[191:188] ^ 3);
  assign w835[31] = |(datain[187:184] ^ 11);
  assign w835[32] = |(datain[183:180] ^ 13);
  assign w835[33] = |(datain[179:176] ^ 10);
  assign w835[34] = |(datain[175:172] ^ 7);
  assign w835[35] = |(datain[171:168] ^ 4);
  assign w835[36] = |(datain[167:164] ^ 0);
  assign w835[37] = |(datain[163:160] ^ 5);
  assign w835[38] = |(datain[159:156] ^ 3);
  assign w835[39] = |(datain[155:152] ^ 0);
  assign w835[40] = |(datain[151:148] ^ 0);
  assign w835[41] = |(datain[147:144] ^ 15);
  assign w835[42] = |(datain[143:140] ^ 4);
  assign w835[43] = |(datain[139:136] ^ 3);
  assign w835[44] = |(datain[135:132] ^ 14);
  assign w835[45] = |(datain[131:128] ^ 11);
  assign w835[46] = |(datain[127:124] ^ 15);
  assign w835[47] = |(datain[123:120] ^ 7);
  assign w835[48] = |(datain[119:116] ^ 9);
  assign w835[49] = |(datain[115:112] ^ 0);
  assign comp[835] = ~(|w835);
  wire [50-1:0] w836;
  assign w836[0] = |(datain[311:308] ^ 0);
  assign w836[1] = |(datain[307:304] ^ 3);
  assign w836[2] = |(datain[303:300] ^ 0);
  assign w836[3] = |(datain[299:296] ^ 1);
  assign w836[4] = |(datain[295:292] ^ 8);
  assign w836[5] = |(datain[291:288] ^ 13);
  assign w836[6] = |(datain[287:284] ^ 9);
  assign w836[7] = |(datain[283:280] ^ 14);
  assign w836[8] = |(datain[279:276] ^ 2);
  assign w836[9] = |(datain[275:272] ^ 0);
  assign w836[10] = |(datain[271:268] ^ 0);
  assign w836[11] = |(datain[267:264] ^ 1);
  assign w836[12] = |(datain[263:260] ^ 8);
  assign w836[13] = |(datain[259:256] ^ 13);
  assign w836[14] = |(datain[255:252] ^ 9);
  assign w836[15] = |(datain[251:248] ^ 6);
  assign w836[16] = |(datain[247:244] ^ 10);
  assign w836[17] = |(datain[243:240] ^ 6);
  assign w836[18] = |(datain[239:236] ^ 0);
  assign w836[19] = |(datain[235:232] ^ 1);
  assign w836[20] = |(datain[231:228] ^ 3);
  assign w836[21] = |(datain[227:224] ^ 14);
  assign w836[22] = |(datain[223:220] ^ 8);
  assign w836[23] = |(datain[219:216] ^ 10);
  assign w836[24] = |(datain[215:212] ^ 8);
  assign w836[25] = |(datain[211:208] ^ 14);
  assign w836[26] = |(datain[207:204] ^ 0);
  assign w836[27] = |(datain[203:200] ^ 3);
  assign w836[28] = |(datain[199:196] ^ 0);
  assign w836[29] = |(datain[195:192] ^ 1);
  assign w836[30] = |(datain[191:188] ^ 3);
  assign w836[31] = |(datain[187:184] ^ 11);
  assign w836[32] = |(datain[183:180] ^ 13);
  assign w836[33] = |(datain[179:176] ^ 10);
  assign w836[34] = |(datain[175:172] ^ 7);
  assign w836[35] = |(datain[171:168] ^ 4);
  assign w836[36] = |(datain[167:164] ^ 0);
  assign w836[37] = |(datain[163:160] ^ 5);
  assign w836[38] = |(datain[159:156] ^ 3);
  assign w836[39] = |(datain[155:152] ^ 0);
  assign w836[40] = |(datain[151:148] ^ 0);
  assign w836[41] = |(datain[147:144] ^ 15);
  assign w836[42] = |(datain[143:140] ^ 4);
  assign w836[43] = |(datain[139:136] ^ 3);
  assign w836[44] = |(datain[135:132] ^ 14);
  assign w836[45] = |(datain[131:128] ^ 11);
  assign w836[46] = |(datain[127:124] ^ 15);
  assign w836[47] = |(datain[123:120] ^ 7);
  assign w836[48] = |(datain[119:116] ^ 9);
  assign w836[49] = |(datain[115:112] ^ 0);
  assign comp[836] = ~(|w836);
  wire [46-1:0] w837;
  assign w837[0] = |(datain[311:308] ^ 8);
  assign w837[1] = |(datain[307:304] ^ 1);
  assign w837[2] = |(datain[303:300] ^ 14);
  assign w837[3] = |(datain[299:296] ^ 13);
  assign w837[4] = |(datain[295:292] ^ 0);
  assign w837[5] = |(datain[291:288] ^ 3);
  assign w837[6] = |(datain[287:284] ^ 0);
  assign w837[7] = |(datain[283:280] ^ 1);
  assign w837[8] = |(datain[279:276] ^ 8);
  assign w837[9] = |(datain[275:272] ^ 13);
  assign w837[10] = |(datain[271:268] ^ 9);
  assign w837[11] = |(datain[267:264] ^ 14);
  assign w837[12] = |(datain[263:260] ^ 2);
  assign w837[13] = |(datain[259:256] ^ 0);
  assign w837[14] = |(datain[255:252] ^ 0);
  assign w837[15] = |(datain[251:248] ^ 1);
  assign w837[16] = |(datain[247:244] ^ 8);
  assign w837[17] = |(datain[243:240] ^ 13);
  assign w837[18] = |(datain[239:236] ^ 9);
  assign w837[19] = |(datain[235:232] ^ 6);
  assign w837[20] = |(datain[231:228] ^ 8);
  assign w837[21] = |(datain[227:224] ^ 11);
  assign w837[22] = |(datain[223:220] ^ 0);
  assign w837[23] = |(datain[219:216] ^ 1);
  assign w837[24] = |(datain[215:212] ^ 3);
  assign w837[25] = |(datain[211:208] ^ 14);
  assign w837[26] = |(datain[207:204] ^ 8);
  assign w837[27] = |(datain[203:200] ^ 10);
  assign w837[28] = |(datain[199:196] ^ 8);
  assign w837[29] = |(datain[195:192] ^ 14);
  assign w837[30] = |(datain[191:188] ^ 0);
  assign w837[31] = |(datain[187:184] ^ 3);
  assign w837[32] = |(datain[183:180] ^ 0);
  assign w837[33] = |(datain[179:176] ^ 1);
  assign w837[34] = |(datain[175:172] ^ 3);
  assign w837[35] = |(datain[171:168] ^ 11);
  assign w837[36] = |(datain[167:164] ^ 13);
  assign w837[37] = |(datain[163:160] ^ 10);
  assign w837[38] = |(datain[159:156] ^ 7);
  assign w837[39] = |(datain[155:152] ^ 4);
  assign w837[40] = |(datain[151:148] ^ 0);
  assign w837[41] = |(datain[147:144] ^ 5);
  assign w837[42] = |(datain[143:140] ^ 3);
  assign w837[43] = |(datain[139:136] ^ 0);
  assign w837[44] = |(datain[135:132] ^ 0);
  assign w837[45] = |(datain[131:128] ^ 15);
  assign comp[837] = ~(|w837);
  wire [62-1:0] w838;
  assign w838[0] = |(datain[311:308] ^ 1);
  assign w838[1] = |(datain[307:304] ^ 4);
  assign w838[2] = |(datain[303:300] ^ 2);
  assign w838[3] = |(datain[299:296] ^ 0);
  assign w838[4] = |(datain[295:292] ^ 1);
  assign w838[5] = |(datain[291:288] ^ 14);
  assign w838[6] = |(datain[287:284] ^ 5);
  assign w838[7] = |(datain[283:280] ^ 7);
  assign w838[8] = |(datain[279:276] ^ 11);
  assign w838[9] = |(datain[275:272] ^ 15);
  assign w838[10] = |(datain[271:268] ^ 5);
  assign w838[11] = |(datain[267:264] ^ 4);
  assign w838[12] = |(datain[263:260] ^ 0);
  assign w838[13] = |(datain[259:256] ^ 0);
  assign w838[14] = |(datain[255:252] ^ 1);
  assign w838[15] = |(datain[251:248] ^ 14);
  assign w838[16] = |(datain[247:244] ^ 5);
  assign w838[17] = |(datain[243:240] ^ 7);
  assign w838[18] = |(datain[239:236] ^ 11);
  assign w838[19] = |(datain[235:232] ^ 8);
  assign w838[20] = |(datain[231:228] ^ 8);
  assign w838[21] = |(datain[227:224] ^ 8);
  assign w838[22] = |(datain[223:220] ^ 1);
  assign w838[23] = |(datain[219:216] ^ 3);
  assign w838[24] = |(datain[215:212] ^ 5);
  assign w838[25] = |(datain[211:208] ^ 0);
  assign w838[26] = |(datain[207:204] ^ 11);
  assign w838[27] = |(datain[203:200] ^ 15);
  assign w838[28] = |(datain[199:196] ^ 9);
  assign w838[29] = |(datain[195:192] ^ 6);
  assign w838[30] = |(datain[191:188] ^ 2);
  assign w838[31] = |(datain[187:184] ^ 0);
  assign w838[32] = |(datain[183:180] ^ 1);
  assign w838[33] = |(datain[179:176] ^ 14);
  assign w838[34] = |(datain[175:172] ^ 5);
  assign w838[35] = |(datain[171:168] ^ 7);
  assign w838[36] = |(datain[167:164] ^ 9);
  assign w838[37] = |(datain[163:160] ^ 10);
  assign w838[38] = |(datain[159:156] ^ 12);
  assign w838[39] = |(datain[155:152] ^ 0);
  assign w838[40] = |(datain[151:148] ^ 0);
  assign w838[41] = |(datain[147:144] ^ 5);
  assign w838[42] = |(datain[143:140] ^ 6);
  assign w838[43] = |(datain[139:136] ^ 1);
  assign w838[44] = |(datain[135:132] ^ 0);
  assign w838[45] = |(datain[131:128] ^ 0);
  assign w838[46] = |(datain[127:124] ^ 9);
  assign w838[47] = |(datain[123:120] ^ 10);
  assign w838[48] = |(datain[119:116] ^ 9);
  assign w838[49] = |(datain[115:112] ^ 1);
  assign w838[50] = |(datain[111:108] ^ 0);
  assign w838[51] = |(datain[107:104] ^ 2);
  assign w838[52] = |(datain[103:100] ^ 6);
  assign w838[53] = |(datain[99:96] ^ 1);
  assign w838[54] = |(datain[95:92] ^ 0);
  assign w838[55] = |(datain[91:88] ^ 0);
  assign w838[56] = |(datain[87:84] ^ 11);
  assign w838[57] = |(datain[83:80] ^ 15);
  assign w838[58] = |(datain[79:76] ^ 1);
  assign w838[59] = |(datain[75:72] ^ 4);
  assign w838[60] = |(datain[71:68] ^ 2);
  assign w838[61] = |(datain[67:64] ^ 0);
  assign comp[838] = ~(|w838);
  wire [30-1:0] w839;
  assign w839[0] = |(datain[311:308] ^ 7);
  assign w839[1] = |(datain[307:304] ^ 15);
  assign w839[2] = |(datain[303:300] ^ 0);
  assign w839[3] = |(datain[299:296] ^ 2);
  assign w839[4] = |(datain[295:292] ^ 11);
  assign w839[5] = |(datain[291:288] ^ 4);
  assign w839[6] = |(datain[287:284] ^ 3);
  assign w839[7] = |(datain[283:280] ^ 15);
  assign w839[8] = |(datain[279:276] ^ 11);
  assign w839[9] = |(datain[275:272] ^ 9);
  assign w839[10] = |(datain[271:268] ^ 0);
  assign w839[11] = |(datain[267:264] ^ 3);
  assign w839[12] = |(datain[263:260] ^ 0);
  assign w839[13] = |(datain[259:256] ^ 0);
  assign w839[14] = |(datain[255:252] ^ 8);
  assign w839[15] = |(datain[251:248] ^ 13);
  assign w839[16] = |(datain[247:244] ^ 9);
  assign w839[17] = |(datain[243:240] ^ 5);
  assign w839[18] = |(datain[239:236] ^ 8);
  assign w839[19] = |(datain[235:232] ^ 1);
  assign w839[20] = |(datain[231:228] ^ 0);
  assign w839[21] = |(datain[227:224] ^ 2);
  assign w839[22] = |(datain[223:220] ^ 12);
  assign w839[23] = |(datain[219:216] ^ 13);
  assign w839[24] = |(datain[215:212] ^ 2);
  assign w839[25] = |(datain[211:208] ^ 1);
  assign w839[26] = |(datain[207:204] ^ 7);
  assign w839[27] = |(datain[203:200] ^ 2);
  assign w839[28] = |(datain[199:196] ^ 3);
  assign w839[29] = |(datain[195:192] ^ 2);
  assign comp[839] = ~(|w839);
  wire [42-1:0] w840;
  assign w840[0] = |(datain[311:308] ^ 12);
  assign w840[1] = |(datain[307:304] ^ 13);
  assign w840[2] = |(datain[303:300] ^ 2);
  assign w840[3] = |(datain[299:296] ^ 1);
  assign w840[4] = |(datain[295:292] ^ 12);
  assign w840[5] = |(datain[291:288] ^ 3);
  assign w840[6] = |(datain[287:284] ^ 8);
  assign w840[7] = |(datain[283:280] ^ 13);
  assign w840[8] = |(datain[279:276] ^ 11);
  assign w840[9] = |(datain[275:272] ^ 5);
  assign w840[10] = |(datain[271:268] ^ 8);
  assign w840[11] = |(datain[267:264] ^ 4);
  assign w840[12] = |(datain[263:260] ^ 0);
  assign w840[13] = |(datain[259:256] ^ 2);
  assign w840[14] = |(datain[255:252] ^ 5);
  assign w840[15] = |(datain[251:248] ^ 7);
  assign w840[16] = |(datain[247:244] ^ 11);
  assign w840[17] = |(datain[243:240] ^ 9);
  assign w840[18] = |(datain[239:236] ^ 3);
  assign w840[19] = |(datain[235:232] ^ 1);
  assign w840[20] = |(datain[231:228] ^ 0);
  assign w840[21] = |(datain[227:224] ^ 0);
  assign w840[22] = |(datain[223:220] ^ 8);
  assign w840[23] = |(datain[219:216] ^ 11);
  assign w840[24] = |(datain[215:212] ^ 15);
  assign w840[25] = |(datain[211:208] ^ 14);
  assign w840[26] = |(datain[207:204] ^ 10);
  assign w840[27] = |(datain[203:200] ^ 12);
  assign w840[28] = |(datain[199:196] ^ 3);
  assign w840[29] = |(datain[195:192] ^ 4);
  assign w840[30] = |(datain[191:188] ^ 8);
  assign w840[31] = |(datain[187:184] ^ 0);
  assign w840[32] = |(datain[183:180] ^ 10);
  assign w840[33] = |(datain[179:176] ^ 10);
  assign w840[34] = |(datain[175:172] ^ 14);
  assign w840[35] = |(datain[171:168] ^ 2);
  assign w840[36] = |(datain[167:164] ^ 15);
  assign w840[37] = |(datain[163:160] ^ 10);
  assign w840[38] = |(datain[159:156] ^ 5);
  assign w840[39] = |(datain[155:152] ^ 15);
  assign w840[40] = |(datain[151:148] ^ 12);
  assign w840[41] = |(datain[147:144] ^ 3);
  assign comp[840] = ~(|w840);
  wire [44-1:0] w841;
  assign w841[0] = |(datain[311:308] ^ 2);
  assign w841[1] = |(datain[307:304] ^ 14);
  assign w841[2] = |(datain[303:300] ^ 8);
  assign w841[3] = |(datain[299:296] ^ 14);
  assign w841[4] = |(datain[295:292] ^ 5);
  assign w841[5] = |(datain[291:288] ^ 5);
  assign w841[6] = |(datain[287:284] ^ 15);
  assign w841[7] = |(datain[283:280] ^ 8);
  assign w841[8] = |(datain[279:276] ^ 2);
  assign w841[9] = |(datain[275:272] ^ 14);
  assign w841[10] = |(datain[271:268] ^ 8);
  assign w841[11] = |(datain[267:264] ^ 11);
  assign w841[12] = |(datain[263:260] ^ 6);
  assign w841[13] = |(datain[259:256] ^ 5);
  assign w841[14] = |(datain[255:252] ^ 15);
  assign w841[15] = |(datain[251:248] ^ 10);
  assign w841[16] = |(datain[247:244] ^ 15);
  assign w841[17] = |(datain[243:240] ^ 11);
  assign w841[18] = |(datain[239:236] ^ 2);
  assign w841[19] = |(datain[235:232] ^ 14);
  assign w841[20] = |(datain[231:228] ^ 15);
  assign w841[21] = |(datain[227:224] ^ 15);
  assign w841[22] = |(datain[223:220] ^ 6);
  assign w841[23] = |(datain[219:216] ^ 13);
  assign w841[24] = |(datain[215:212] ^ 15);
  assign w841[25] = |(datain[211:208] ^ 12);
  assign w841[26] = |(datain[207:204] ^ 9);
  assign w841[27] = |(datain[203:200] ^ 12);
  assign w841[28] = |(datain[199:196] ^ 8);
  assign w841[29] = |(datain[195:192] ^ 0);
  assign w841[30] = |(datain[191:188] ^ 15);
  assign w841[31] = |(datain[187:184] ^ 12);
  assign w841[32] = |(datain[183:180] ^ 15);
  assign w841[33] = |(datain[179:176] ^ 0);
  assign w841[34] = |(datain[175:172] ^ 7);
  assign w841[35] = |(datain[171:168] ^ 5);
  assign w841[36] = |(datain[167:164] ^ 0);
  assign w841[37] = |(datain[163:160] ^ 4);
  assign w841[38] = |(datain[159:156] ^ 11);
  assign w841[39] = |(datain[155:152] ^ 4);
  assign w841[40] = |(datain[151:148] ^ 1);
  assign w841[41] = |(datain[147:144] ^ 9);
  assign w841[42] = |(datain[143:140] ^ 9);
  assign w841[43] = |(datain[139:136] ^ 13);
  assign comp[841] = ~(|w841);
  wire [32-1:0] w842;
  assign w842[0] = |(datain[311:308] ^ 11);
  assign w842[1] = |(datain[307:304] ^ 4);
  assign w842[2] = |(datain[303:300] ^ 15);
  assign w842[3] = |(datain[299:296] ^ 0);
  assign w842[4] = |(datain[295:292] ^ 12);
  assign w842[5] = |(datain[291:288] ^ 13);
  assign w842[6] = |(datain[287:284] ^ 1);
  assign w842[7] = |(datain[283:280] ^ 3);
  assign w842[8] = |(datain[279:276] ^ 8);
  assign w842[9] = |(datain[275:272] ^ 0);
  assign w842[10] = |(datain[271:268] ^ 15);
  assign w842[11] = |(datain[267:264] ^ 12);
  assign w842[12] = |(datain[263:260] ^ 1);
  assign w842[13] = |(datain[259:256] ^ 9);
  assign w842[14] = |(datain[255:252] ^ 7);
  assign w842[15] = |(datain[251:248] ^ 4);
  assign w842[16] = |(datain[247:244] ^ 1);
  assign w842[17] = |(datain[243:240] ^ 0);
  assign w842[18] = |(datain[239:236] ^ 8);
  assign w842[19] = |(datain[235:232] ^ 12);
  assign w842[20] = |(datain[231:228] ^ 13);
  assign w842[21] = |(datain[227:224] ^ 8);
  assign w842[22] = |(datain[223:220] ^ 4);
  assign w842[23] = |(datain[219:216] ^ 8);
  assign w842[24] = |(datain[215:212] ^ 8);
  assign w842[25] = |(datain[211:208] ^ 14);
  assign w842[26] = |(datain[207:204] ^ 13);
  assign w842[27] = |(datain[203:200] ^ 8);
  assign w842[28] = |(datain[199:196] ^ 2);
  assign w842[29] = |(datain[195:192] ^ 9);
  assign w842[30] = |(datain[191:188] ^ 1);
  assign w842[31] = |(datain[187:184] ^ 6);
  assign comp[842] = ~(|w842);
  wire [48-1:0] w843;
  assign w843[0] = |(datain[311:308] ^ 5);
  assign w843[1] = |(datain[307:304] ^ 1);
  assign w843[2] = |(datain[303:300] ^ 0);
  assign w843[3] = |(datain[299:296] ^ 15);
  assign w843[4] = |(datain[295:292] ^ 8);
  assign w843[5] = |(datain[291:288] ^ 14);
  assign w843[6] = |(datain[287:284] ^ 13);
  assign w843[7] = |(datain[283:280] ^ 10);
  assign w843[8] = |(datain[279:276] ^ 11);
  assign w843[9] = |(datain[275:272] ^ 14);
  assign w843[10] = |(datain[271:268] ^ 1);
  assign w843[11] = |(datain[267:264] ^ 11);
  assign w843[12] = |(datain[263:260] ^ 0);
  assign w843[13] = |(datain[259:256] ^ 0);
  assign w843[14] = |(datain[255:252] ^ 8);
  assign w843[15] = |(datain[251:248] ^ 0);
  assign w843[16] = |(datain[247:244] ^ 0);
  assign w843[17] = |(datain[243:240] ^ 4);
  assign w843[18] = |(datain[239:236] ^ 14);
  assign w843[19] = |(datain[235:232] ^ 7);
  assign w843[20] = |(datain[231:228] ^ 8);
  assign w843[21] = |(datain[227:224] ^ 0);
  assign w843[22] = |(datain[223:220] ^ 2);
  assign w843[23] = |(datain[219:216] ^ 14);
  assign w843[24] = |(datain[215:212] ^ 0);
  assign w843[25] = |(datain[211:208] ^ 12);
  assign w843[26] = |(datain[207:204] ^ 0);
  assign w843[27] = |(datain[203:200] ^ 0);
  assign w843[28] = |(datain[199:196] ^ 15);
  assign w843[29] = |(datain[195:192] ^ 1);
  assign w843[30] = |(datain[191:188] ^ 8);
  assign w843[31] = |(datain[187:184] ^ 3);
  assign w843[32] = |(datain[183:180] ^ 12);
  assign w843[33] = |(datain[179:176] ^ 6);
  assign w843[34] = |(datain[175:172] ^ 0);
  assign w843[35] = |(datain[171:168] ^ 1);
  assign w843[36] = |(datain[167:164] ^ 8);
  assign w843[37] = |(datain[163:160] ^ 1);
  assign w843[38] = |(datain[159:156] ^ 15);
  assign w843[39] = |(datain[155:152] ^ 14);
  assign w843[40] = |(datain[151:148] ^ 5);
  assign w843[41] = |(datain[147:144] ^ 7);
  assign w843[42] = |(datain[143:140] ^ 0);
  assign w843[43] = |(datain[139:136] ^ 8);
  assign w843[44] = |(datain[135:132] ^ 7);
  assign w843[45] = |(datain[131:128] ^ 6);
  assign w843[46] = |(datain[127:124] ^ 14);
  assign w843[47] = |(datain[123:120] ^ 15);
  assign comp[843] = ~(|w843);
  wire [30-1:0] w844;
  assign w844[0] = |(datain[311:308] ^ 8);
  assign w844[1] = |(datain[307:304] ^ 0);
  assign w844[2] = |(datain[303:300] ^ 15);
  assign w844[3] = |(datain[299:296] ^ 12);
  assign w844[4] = |(datain[295:292] ^ 4);
  assign w844[5] = |(datain[291:288] ^ 11);
  assign w844[6] = |(datain[287:284] ^ 7);
  assign w844[7] = |(datain[283:280] ^ 4);
  assign w844[8] = |(datain[279:276] ^ 1);
  assign w844[9] = |(datain[275:272] ^ 2);
  assign w844[10] = |(datain[271:268] ^ 3);
  assign w844[11] = |(datain[267:264] ^ 13);
  assign w844[12] = |(datain[263:260] ^ 0);
  assign w844[13] = |(datain[259:256] ^ 0);
  assign w844[14] = |(datain[255:252] ^ 3);
  assign w844[15] = |(datain[251:248] ^ 13);
  assign w844[16] = |(datain[247:244] ^ 7);
  assign w844[17] = |(datain[243:240] ^ 4);
  assign w844[18] = |(datain[239:236] ^ 0);
  assign w844[19] = |(datain[235:232] ^ 13);
  assign w844[20] = |(datain[231:228] ^ 3);
  assign w844[21] = |(datain[227:224] ^ 13);
  assign w844[22] = |(datain[223:220] ^ 0);
  assign w844[23] = |(datain[219:216] ^ 0);
  assign w844[24] = |(datain[215:212] ^ 6);
  assign w844[25] = |(datain[211:208] ^ 12);
  assign w844[26] = |(datain[207:204] ^ 7);
  assign w844[27] = |(datain[203:200] ^ 5);
  assign w844[28] = |(datain[199:196] ^ 0);
  assign w844[29] = |(datain[195:192] ^ 5);
  assign comp[844] = ~(|w844);
  wire [42-1:0] w845;
  assign w845[0] = |(datain[311:308] ^ 0);
  assign w845[1] = |(datain[307:304] ^ 14);
  assign w845[2] = |(datain[303:300] ^ 1);
  assign w845[3] = |(datain[299:296] ^ 15);
  assign w845[4] = |(datain[295:292] ^ 14);
  assign w845[5] = |(datain[291:288] ^ 8);
  assign w845[6] = |(datain[287:284] ^ 0);
  assign w845[7] = |(datain[283:280] ^ 0);
  assign w845[8] = |(datain[279:276] ^ 0);
  assign w845[9] = |(datain[275:272] ^ 0);
  assign w845[10] = |(datain[271:268] ^ 5);
  assign w845[11] = |(datain[267:264] ^ 14);
  assign w845[12] = |(datain[263:260] ^ 11);
  assign w845[13] = |(datain[259:256] ^ 9);
  assign w845[14] = |(datain[255:252] ^ 14);
  assign w845[15] = |(datain[251:248] ^ 0);
  assign w845[16] = |(datain[247:244] ^ 0);
  assign w845[17] = |(datain[243:240] ^ 1);
  assign w845[18] = |(datain[239:236] ^ 8);
  assign w845[19] = |(datain[235:232] ^ 3);
  assign w845[20] = |(datain[231:228] ^ 12);
  assign w845[21] = |(datain[227:224] ^ 6);
  assign w845[22] = |(datain[223:220] ^ 1);
  assign w845[23] = |(datain[219:216] ^ 1);
  assign w845[24] = |(datain[215:212] ^ 9);
  assign w845[25] = |(datain[211:208] ^ 0);
  assign w845[26] = |(datain[207:204] ^ 8);
  assign w845[27] = |(datain[203:200] ^ 1);
  assign w845[28] = |(datain[199:196] ^ 3);
  assign w845[29] = |(datain[195:192] ^ 4);
  assign w845[30] = |(datain[191:188] ^ 1);
  assign w845[31] = |(datain[187:184] ^ 1);
  assign w845[32] = |(datain[183:180] ^ 2);
  assign w845[33] = |(datain[179:176] ^ 3);
  assign w845[34] = |(datain[175:172] ^ 4);
  assign w845[35] = |(datain[171:168] ^ 6);
  assign w845[36] = |(datain[167:164] ^ 4);
  assign w845[37] = |(datain[163:160] ^ 6);
  assign w845[38] = |(datain[159:156] ^ 14);
  assign w845[39] = |(datain[155:152] ^ 2);
  assign w845[40] = |(datain[151:148] ^ 15);
  assign w845[41] = |(datain[147:144] ^ 8);
  assign comp[845] = ~(|w845);
  wire [34-1:0] w846;
  assign w846[0] = |(datain[311:308] ^ 5);
  assign w846[1] = |(datain[307:304] ^ 11);
  assign w846[2] = |(datain[303:300] ^ 8);
  assign w846[3] = |(datain[299:296] ^ 3);
  assign w846[4] = |(datain[295:292] ^ 12);
  assign w846[5] = |(datain[291:288] ^ 3);
  assign w846[6] = |(datain[287:284] ^ 1);
  assign w846[7] = |(datain[283:280] ^ 1);
  assign w846[8] = |(datain[279:276] ^ 11);
  assign w846[9] = |(datain[275:272] ^ 9);
  assign w846[10] = |(datain[271:268] ^ 10);
  assign w846[11] = |(datain[267:264] ^ 8);
  assign w846[12] = |(datain[263:260] ^ 0);
  assign w846[13] = |(datain[259:256] ^ 1);
  assign w846[14] = |(datain[255:252] ^ 0);
  assign w846[15] = |(datain[251:248] ^ 14);
  assign w846[16] = |(datain[247:244] ^ 1);
  assign w846[17] = |(datain[243:240] ^ 15);
  assign w846[18] = |(datain[239:236] ^ 8);
  assign w846[19] = |(datain[235:232] ^ 1);
  assign w846[20] = |(datain[231:228] ^ 3);
  assign w846[21] = |(datain[227:224] ^ 7);
  assign w846[22] = |(datain[223:220] ^ 2);
  assign w846[23] = |(datain[219:216] ^ 0);
  assign w846[24] = |(datain[215:212] ^ 2);
  assign w846[25] = |(datain[211:208] ^ 9);
  assign w846[26] = |(datain[207:204] ^ 4);
  assign w846[27] = |(datain[203:200] ^ 3);
  assign w846[28] = |(datain[199:196] ^ 4);
  assign w846[29] = |(datain[195:192] ^ 3);
  assign w846[30] = |(datain[191:188] ^ 14);
  assign w846[31] = |(datain[187:184] ^ 2);
  assign w846[32] = |(datain[183:180] ^ 15);
  assign w846[33] = |(datain[179:176] ^ 8);
  assign comp[846] = ~(|w846);
  wire [40-1:0] w847;
  assign w847[0] = |(datain[311:308] ^ 14);
  assign w847[1] = |(datain[307:304] ^ 8);
  assign w847[2] = |(datain[303:300] ^ 0);
  assign w847[3] = |(datain[299:296] ^ 0);
  assign w847[4] = |(datain[295:292] ^ 0);
  assign w847[5] = |(datain[291:288] ^ 0);
  assign w847[6] = |(datain[287:284] ^ 5);
  assign w847[7] = |(datain[283:280] ^ 11);
  assign w847[8] = |(datain[279:276] ^ 11);
  assign w847[9] = |(datain[275:272] ^ 9);
  assign w847[10] = |(datain[271:268] ^ 10);
  assign w847[11] = |(datain[267:264] ^ 8);
  assign w847[12] = |(datain[263:260] ^ 0);
  assign w847[13] = |(datain[259:256] ^ 1);
  assign w847[14] = |(datain[255:252] ^ 0);
  assign w847[15] = |(datain[251:248] ^ 14);
  assign w847[16] = |(datain[247:244] ^ 1);
  assign w847[17] = |(datain[243:240] ^ 15);
  assign w847[18] = |(datain[239:236] ^ 8);
  assign w847[19] = |(datain[235:232] ^ 3);
  assign w847[20] = |(datain[231:228] ^ 12);
  assign w847[21] = |(datain[227:224] ^ 3);
  assign w847[22] = |(datain[223:220] ^ 1);
  assign w847[23] = |(datain[219:216] ^ 1);
  assign w847[24] = |(datain[215:212] ^ 8);
  assign w847[25] = |(datain[211:208] ^ 1);
  assign w847[26] = |(datain[207:204] ^ 3);
  assign w847[27] = |(datain[203:200] ^ 7);
  assign w847[28] = |(datain[199:196] ^ 9);
  assign w847[29] = |(datain[195:192] ^ 3);
  assign w847[30] = |(datain[191:188] ^ 1);
  assign w847[31] = |(datain[187:184] ^ 9);
  assign w847[32] = |(datain[183:180] ^ 4);
  assign w847[33] = |(datain[179:176] ^ 3);
  assign w847[34] = |(datain[175:172] ^ 4);
  assign w847[35] = |(datain[171:168] ^ 3);
  assign w847[36] = |(datain[167:164] ^ 14);
  assign w847[37] = |(datain[163:160] ^ 2);
  assign w847[38] = |(datain[159:156] ^ 15);
  assign w847[39] = |(datain[155:152] ^ 8);
  assign comp[847] = ~(|w847);
  wire [70-1:0] w848;
  assign w848[0] = |(datain[311:308] ^ 5);
  assign w848[1] = |(datain[307:304] ^ 10);
  assign w848[2] = |(datain[303:300] ^ 0);
  assign w848[3] = |(datain[299:296] ^ 14);
  assign w848[4] = |(datain[295:292] ^ 1);
  assign w848[5] = |(datain[291:288] ^ 15);
  assign w848[6] = |(datain[287:284] ^ 11);
  assign w848[7] = |(datain[283:280] ^ 8);
  assign w848[8] = |(datain[279:276] ^ 15);
  assign w848[9] = |(datain[275:272] ^ 15);
  assign w848[10] = |(datain[271:268] ^ 2);
  assign w848[11] = |(datain[267:264] ^ 5);
  assign w848[12] = |(datain[263:260] ^ 8);
  assign w848[13] = |(datain[259:256] ^ 3);
  assign w848[14] = |(datain[255:252] ^ 12);
  assign w848[15] = |(datain[251:248] ^ 2);
  assign w848[16] = |(datain[247:244] ^ 1);
  assign w848[17] = |(datain[243:240] ^ 1);
  assign w848[18] = |(datain[239:236] ^ 9);
  assign w848[19] = |(datain[235:232] ^ 0);
  assign w848[20] = |(datain[231:228] ^ 12);
  assign w848[21] = |(datain[227:224] ^ 13);
  assign w848[22] = |(datain[223:220] ^ 2);
  assign w848[23] = |(datain[219:216] ^ 1);
  assign w848[24] = |(datain[215:212] ^ 12);
  assign w848[25] = |(datain[211:208] ^ 13);
  assign w848[26] = |(datain[207:204] ^ 15);
  assign w848[27] = |(datain[203:200] ^ 15);
  assign w848[28] = |(datain[199:196] ^ 14);
  assign w848[29] = |(datain[195:192] ^ 11);
  assign w848[30] = |(datain[191:188] ^ 1);
  assign w848[31] = |(datain[187:184] ^ 3);
  assign w848[32] = |(datain[183:180] ^ 9);
  assign w848[33] = |(datain[179:176] ^ 0);
  assign w848[34] = |(datain[175:172] ^ 11);
  assign w848[35] = |(datain[171:168] ^ 9);
  assign w848[36] = |(datain[167:164] ^ 14);
  assign w848[37] = |(datain[163:160] ^ 0);
  assign w848[38] = |(datain[159:156] ^ 0);
  assign w848[39] = |(datain[155:152] ^ 1);
  assign w848[40] = |(datain[151:148] ^ 8);
  assign w848[41] = |(datain[147:144] ^ 11);
  assign w848[42] = |(datain[143:140] ^ 15);
  assign w848[43] = |(datain[139:136] ^ 2);
  assign w848[44] = |(datain[135:132] ^ 8);
  assign w848[45] = |(datain[131:128] ^ 3);
  assign w848[46] = |(datain[127:124] ^ 12);
  assign w848[47] = |(datain[123:120] ^ 6);
  assign w848[48] = |(datain[119:116] ^ 1);
  assign w848[49] = |(datain[115:112] ^ 2);
  assign w848[50] = |(datain[111:108] ^ 9);
  assign w848[51] = |(datain[107:104] ^ 0);
  assign w848[52] = |(datain[103:100] ^ 8);
  assign w848[53] = |(datain[99:96] ^ 1);
  assign w848[54] = |(datain[95:92] ^ 3);
  assign w848[55] = |(datain[91:88] ^ 4);
  assign w848[56] = |(datain[87:84] ^ 9);
  assign w848[57] = |(datain[83:80] ^ 3);
  assign w848[58] = |(datain[79:76] ^ 1);
  assign w848[59] = |(datain[75:72] ^ 9);
  assign w848[60] = |(datain[71:68] ^ 4);
  assign w848[61] = |(datain[67:64] ^ 6);
  assign w848[62] = |(datain[63:60] ^ 4);
  assign w848[63] = |(datain[59:56] ^ 6);
  assign w848[64] = |(datain[55:52] ^ 14);
  assign w848[65] = |(datain[51:48] ^ 2);
  assign w848[66] = |(datain[47:44] ^ 15);
  assign w848[67] = |(datain[43:40] ^ 8);
  assign w848[68] = |(datain[39:36] ^ 12);
  assign w848[69] = |(datain[35:32] ^ 15);
  assign comp[848] = ~(|w848);
  wire [38-1:0] w849;
  assign w849[0] = |(datain[311:308] ^ 0);
  assign w849[1] = |(datain[307:304] ^ 2);
  assign w849[2] = |(datain[303:300] ^ 0);
  assign w849[3] = |(datain[299:296] ^ 0);
  assign w849[4] = |(datain[295:292] ^ 0);
  assign w849[5] = |(datain[291:288] ^ 0);
  assign w849[6] = |(datain[287:284] ^ 6);
  assign w849[7] = |(datain[283:280] ^ 0);
  assign w849[8] = |(datain[279:276] ^ 15);
  assign w849[9] = |(datain[275:272] ^ 10);
  assign w849[10] = |(datain[271:268] ^ 11);
  assign w849[11] = |(datain[267:264] ^ 9);
  assign w849[12] = |(datain[263:260] ^ 8);
  assign w849[13] = |(datain[259:256] ^ 12);
  assign w849[14] = |(datain[255:252] ^ 0);
  assign w849[15] = |(datain[251:248] ^ 5);
  assign w849[16] = |(datain[247:244] ^ 5);
  assign w849[17] = |(datain[243:240] ^ 14);
  assign w849[18] = |(datain[239:236] ^ 8);
  assign w849[19] = |(datain[235:232] ^ 3);
  assign w849[20] = |(datain[231:228] ^ 12);
  assign w849[21] = |(datain[227:224] ^ 6);
  assign w849[22] = |(datain[223:220] ^ 1);
  assign w849[23] = |(datain[219:216] ^ 1);
  assign w849[24] = |(datain[215:212] ^ 8);
  assign w849[25] = |(datain[211:208] ^ 1);
  assign w849[26] = |(datain[207:204] ^ 2);
  assign w849[27] = |(datain[203:200] ^ 12);
  assign w849[28] = |(datain[199:196] ^ 3);
  assign w849[29] = |(datain[195:192] ^ 0);
  assign w849[30] = |(datain[191:188] ^ 0);
  assign w849[31] = |(datain[187:184] ^ 12);
  assign w849[32] = |(datain[183:180] ^ 4);
  assign w849[33] = |(datain[179:176] ^ 6);
  assign w849[34] = |(datain[175:172] ^ 14);
  assign w849[35] = |(datain[171:168] ^ 2);
  assign w849[36] = |(datain[167:164] ^ 15);
  assign w849[37] = |(datain[163:160] ^ 9);
  assign comp[849] = ~(|w849);
  wire [50-1:0] w850;
  assign w850[0] = |(datain[311:308] ^ 15);
  assign w850[1] = |(datain[307:304] ^ 10);
  assign w850[2] = |(datain[303:300] ^ 11);
  assign w850[3] = |(datain[299:296] ^ 15);
  assign w850[4] = |(datain[295:292] ^ 1);
  assign w850[5] = |(datain[291:288] ^ 9);
  assign w850[6] = |(datain[287:284] ^ 0);
  assign w850[7] = |(datain[283:280] ^ 1);
  assign w850[8] = |(datain[279:276] ^ 8);
  assign w850[9] = |(datain[275:272] ^ 11);
  assign w850[10] = |(datain[271:268] ^ 15);
  assign w850[11] = |(datain[267:264] ^ 7);
  assign w850[12] = |(datain[263:260] ^ 10);
  assign w850[13] = |(datain[259:256] ^ 13);
  assign w850[14] = |(datain[255:252] ^ 3);
  assign w850[15] = |(datain[251:248] ^ 5);
  assign w850[16] = |(datain[247:244] ^ 5);
  assign w850[17] = |(datain[243:240] ^ 13);
  assign w850[18] = |(datain[239:236] ^ 11);
  assign w850[19] = |(datain[235:232] ^ 0);
  assign w850[20] = |(datain[231:228] ^ 10);
  assign w850[21] = |(datain[227:224] ^ 11);
  assign w850[22] = |(datain[223:220] ^ 10);
  assign w850[23] = |(datain[219:216] ^ 13);
  assign w850[24] = |(datain[215:212] ^ 11);
  assign w850[25] = |(datain[211:208] ^ 1);
  assign w850[26] = |(datain[207:204] ^ 0);
  assign w850[27] = |(datain[203:200] ^ 3);
  assign w850[28] = |(datain[199:196] ^ 13);
  assign w850[29] = |(datain[195:192] ^ 2);
  assign w850[30] = |(datain[191:188] ^ 12);
  assign w850[31] = |(datain[187:184] ^ 8);
  assign w850[32] = |(datain[183:180] ^ 10);
  assign w850[33] = |(datain[179:176] ^ 11);
  assign w850[34] = |(datain[175:172] ^ 14);
  assign w850[35] = |(datain[171:168] ^ 11);
  assign w850[36] = |(datain[167:164] ^ 0);
  assign w850[37] = |(datain[163:160] ^ 0);
  assign w850[38] = |(datain[159:156] ^ 11);
  assign w850[39] = |(datain[155:152] ^ 15);
  assign w850[40] = |(datain[151:148] ^ 2);
  assign w850[41] = |(datain[147:144] ^ 5);
  assign w850[42] = |(datain[143:140] ^ 0);
  assign w850[43] = |(datain[139:136] ^ 1);
  assign w850[44] = |(datain[135:132] ^ 8);
  assign w850[45] = |(datain[131:128] ^ 11);
  assign w850[46] = |(datain[127:124] ^ 14);
  assign w850[47] = |(datain[123:120] ^ 7);
  assign w850[48] = |(datain[119:116] ^ 5);
  assign w850[49] = |(datain[115:112] ^ 8);
  assign comp[850] = ~(|w850);
  wire [50-1:0] w851;
  assign w851[0] = |(datain[311:308] ^ 0);
  assign w851[1] = |(datain[307:304] ^ 1);
  assign w851[2] = |(datain[303:300] ^ 8);
  assign w851[3] = |(datain[299:296] ^ 11);
  assign w851[4] = |(datain[295:292] ^ 15);
  assign w851[5] = |(datain[291:288] ^ 7);
  assign w851[6] = |(datain[287:284] ^ 10);
  assign w851[7] = |(datain[283:280] ^ 13);
  assign w851[8] = |(datain[279:276] ^ 3);
  assign w851[9] = |(datain[275:272] ^ 5);
  assign w851[10] = |(datain[271:268] ^ 5);
  assign w851[11] = |(datain[267:264] ^ 13);
  assign w851[12] = |(datain[263:260] ^ 11);
  assign w851[13] = |(datain[259:256] ^ 0);
  assign w851[14] = |(datain[255:252] ^ 10);
  assign w851[15] = |(datain[251:248] ^ 11);
  assign w851[16] = |(datain[247:244] ^ 10);
  assign w851[17] = |(datain[243:240] ^ 13);
  assign w851[18] = |(datain[239:236] ^ 11);
  assign w851[19] = |(datain[235:232] ^ 1);
  assign w851[20] = |(datain[231:228] ^ 0);
  assign w851[21] = |(datain[227:224] ^ 3);
  assign w851[22] = |(datain[223:220] ^ 13);
  assign w851[23] = |(datain[219:216] ^ 2);
  assign w851[24] = |(datain[215:212] ^ 12);
  assign w851[25] = |(datain[211:208] ^ 8);
  assign w851[26] = |(datain[207:204] ^ 10);
  assign w851[27] = |(datain[203:200] ^ 11);
  assign w851[28] = |(datain[199:196] ^ 14);
  assign w851[29] = |(datain[195:192] ^ 11);
  assign w851[30] = |(datain[191:188] ^ 0);
  assign w851[31] = |(datain[187:184] ^ 0);
  assign w851[32] = |(datain[183:180] ^ 11);
  assign w851[33] = |(datain[179:176] ^ 15);
  assign w851[34] = |(datain[175:172] ^ 2);
  assign w851[35] = |(datain[171:168] ^ 5);
  assign w851[36] = |(datain[167:164] ^ 0);
  assign w851[37] = |(datain[163:160] ^ 1);
  assign w851[38] = |(datain[159:156] ^ 8);
  assign w851[39] = |(datain[155:152] ^ 11);
  assign w851[40] = |(datain[151:148] ^ 14);
  assign w851[41] = |(datain[147:144] ^ 7);
  assign w851[42] = |(datain[143:140] ^ 5);
  assign w851[43] = |(datain[139:136] ^ 8);
  assign w851[44] = |(datain[135:132] ^ 12);
  assign w851[45] = |(datain[131:128] ^ 13);
  assign w851[46] = |(datain[127:124] ^ 2);
  assign w851[47] = |(datain[123:120] ^ 0);
  assign w851[48] = |(datain[119:116] ^ 10);
  assign w851[49] = |(datain[115:112] ^ 9);
  assign comp[851] = ~(|w851);
  wire [44-1:0] w852;
  assign w852[0] = |(datain[311:308] ^ 14);
  assign w852[1] = |(datain[307:304] ^ 8);
  assign w852[2] = |(datain[303:300] ^ 13);
  assign w852[3] = |(datain[299:296] ^ 12);
  assign w852[4] = |(datain[295:292] ^ 0);
  assign w852[5] = |(datain[291:288] ^ 5);
  assign w852[6] = |(datain[287:284] ^ 2);
  assign w852[7] = |(datain[283:280] ^ 14);
  assign w852[8] = |(datain[279:276] ^ 12);
  assign w852[9] = |(datain[275:272] ^ 7);
  assign w852[10] = |(datain[271:268] ^ 0);
  assign w852[11] = |(datain[267:264] ^ 6);
  assign w852[12] = |(datain[263:260] ^ 13);
  assign w852[13] = |(datain[259:256] ^ 14);
  assign w852[14] = |(datain[255:252] ^ 0);
  assign w852[15] = |(datain[251:248] ^ 8);
  assign w852[16] = |(datain[247:244] ^ 3);
  assign w852[17] = |(datain[243:240] ^ 3);
  assign w852[18] = |(datain[239:236] ^ 0);
  assign w852[19] = |(datain[235:232] ^ 0);
  assign w852[20] = |(datain[231:228] ^ 9);
  assign w852[21] = |(datain[227:224] ^ 12);
  assign w852[22] = |(datain[223:220] ^ 5);
  assign w852[23] = |(datain[219:216] ^ 8);
  assign w852[24] = |(datain[215:212] ^ 0);
  assign w852[25] = |(datain[211:208] ^ 13);
  assign w852[26] = |(datain[207:204] ^ 0);
  assign w852[27] = |(datain[203:200] ^ 0);
  assign w852[28] = |(datain[199:196] ^ 0);
  assign w852[29] = |(datain[195:192] ^ 3);
  assign w852[30] = |(datain[191:188] ^ 5);
  assign w852[31] = |(datain[187:184] ^ 0);
  assign w852[32] = |(datain[183:180] ^ 9);
  assign w852[33] = |(datain[179:176] ^ 13);
  assign w852[34] = |(datain[175:172] ^ 9);
  assign w852[35] = |(datain[171:168] ^ 0);
  assign w852[36] = |(datain[167:164] ^ 9);
  assign w852[37] = |(datain[163:160] ^ 0);
  assign w852[38] = |(datain[159:156] ^ 9);
  assign w852[39] = |(datain[155:152] ^ 0);
  assign w852[40] = |(datain[151:148] ^ 9);
  assign w852[41] = |(datain[147:144] ^ 0);
  assign w852[42] = |(datain[143:140] ^ 9);
  assign w852[43] = |(datain[139:136] ^ 0);
  assign comp[852] = ~(|w852);
  wire [48-1:0] w853;
  assign w853[0] = |(datain[311:308] ^ 11);
  assign w853[1] = |(datain[307:304] ^ 9);
  assign w853[2] = |(datain[303:300] ^ 0);
  assign w853[3] = |(datain[299:296] ^ 0);
  assign w853[4] = |(datain[295:292] ^ 0);
  assign w853[5] = |(datain[291:288] ^ 4);
  assign w853[6] = |(datain[287:284] ^ 5);
  assign w853[7] = |(datain[283:280] ^ 1);
  assign w853[8] = |(datain[279:276] ^ 5);
  assign w853[9] = |(datain[275:272] ^ 6);
  assign w853[10] = |(datain[271:268] ^ 15);
  assign w853[11] = |(datain[267:264] ^ 11);
  assign w853[12] = |(datain[263:260] ^ 15);
  assign w853[13] = |(datain[259:256] ^ 12);
  assign w853[14] = |(datain[255:252] ^ 15);
  assign w853[15] = |(datain[251:248] ^ 3);
  assign w853[16] = |(datain[247:244] ^ 10);
  assign w853[17] = |(datain[243:240] ^ 5);
  assign w853[18] = |(datain[239:236] ^ 5);
  assign w853[19] = |(datain[235:232] ^ 14);
  assign w853[20] = |(datain[231:228] ^ 5);
  assign w853[21] = |(datain[227:224] ^ 9);
  assign w853[22] = |(datain[223:220] ^ 15);
  assign w853[23] = |(datain[219:216] ^ 12);
  assign w853[24] = |(datain[215:212] ^ 15);
  assign w853[25] = |(datain[211:208] ^ 3);
  assign w853[26] = |(datain[207:204] ^ 10);
  assign w853[27] = |(datain[203:200] ^ 5);
  assign w853[28] = |(datain[199:196] ^ 8);
  assign w853[29] = |(datain[195:192] ^ 11);
  assign w853[30] = |(datain[191:188] ^ 4);
  assign w853[31] = |(datain[187:184] ^ 4);
  assign w853[32] = |(datain[183:180] ^ 15);
  assign w853[33] = |(datain[179:176] ^ 14);
  assign w853[34] = |(datain[175:172] ^ 11);
  assign w853[35] = |(datain[171:168] ^ 9);
  assign w853[36] = |(datain[167:164] ^ 9);
  assign w853[37] = |(datain[163:160] ^ 14);
  assign w853[38] = |(datain[159:156] ^ 0);
  assign w853[39] = |(datain[155:152] ^ 3);
  assign w853[40] = |(datain[151:148] ^ 11);
  assign w853[41] = |(datain[147:144] ^ 11);
  assign w853[42] = |(datain[143:140] ^ 0);
  assign w853[43] = |(datain[139:136] ^ 4);
  assign w853[44] = |(datain[135:132] ^ 0);
  assign w853[45] = |(datain[131:128] ^ 0);
  assign w853[46] = |(datain[127:124] ^ 0);
  assign w853[47] = |(datain[123:120] ^ 6);
  assign comp[853] = ~(|w853);
  wire [76-1:0] w854;
  assign w854[0] = |(datain[311:308] ^ 0);
  assign w854[1] = |(datain[307:304] ^ 1);
  assign w854[2] = |(datain[303:300] ^ 14);
  assign w854[3] = |(datain[299:296] ^ 8);
  assign w854[4] = |(datain[295:292] ^ 0);
  assign w854[5] = |(datain[291:288] ^ 9);
  assign w854[6] = |(datain[287:284] ^ 0);
  assign w854[7] = |(datain[283:280] ^ 0);
  assign w854[8] = |(datain[279:276] ^ 0);
  assign w854[9] = |(datain[275:272] ^ 7);
  assign w854[10] = |(datain[271:268] ^ 14);
  assign w854[11] = |(datain[267:264] ^ 8);
  assign w854[12] = |(datain[263:260] ^ 0);
  assign w854[13] = |(datain[259:256] ^ 14);
  assign w854[14] = |(datain[255:252] ^ 0);
  assign w854[15] = |(datain[251:248] ^ 0);
  assign w854[16] = |(datain[247:244] ^ 14);
  assign w854[17] = |(datain[243:240] ^ 10);
  assign w854[18] = |(datain[239:236] ^ 0);
  assign w854[19] = |(datain[235:232] ^ 0);
  assign w854[20] = |(datain[231:228] ^ 0);
  assign w854[21] = |(datain[227:224] ^ 0);
  assign w854[22] = |(datain[223:220] ^ 15);
  assign w854[23] = |(datain[219:216] ^ 15);
  assign w854[24] = |(datain[215:212] ^ 15);
  assign w854[25] = |(datain[211:208] ^ 15);
  assign w854[26] = |(datain[207:204] ^ 10);
  assign w854[27] = |(datain[203:200] ^ 5);
  assign w854[28] = |(datain[199:196] ^ 10);
  assign w854[29] = |(datain[195:192] ^ 5);
  assign w854[30] = |(datain[191:188] ^ 8);
  assign w854[31] = |(datain[187:184] ^ 9);
  assign w854[32] = |(datain[183:180] ^ 4);
  assign w854[33] = |(datain[179:176] ^ 4);
  assign w854[34] = |(datain[175:172] ^ 15);
  assign w854[35] = |(datain[171:168] ^ 12);
  assign w854[36] = |(datain[167:164] ^ 8);
  assign w854[37] = |(datain[163:160] ^ 12);
  assign w854[38] = |(datain[159:156] ^ 4);
  assign w854[39] = |(datain[155:152] ^ 4);
  assign w854[40] = |(datain[151:148] ^ 15);
  assign w854[41] = |(datain[147:144] ^ 14);
  assign w854[42] = |(datain[143:140] ^ 12);
  assign w854[43] = |(datain[139:136] ^ 3);
  assign w854[44] = |(datain[135:132] ^ 0);
  assign w854[45] = |(datain[131:128] ^ 14);
  assign w854[46] = |(datain[127:124] ^ 1);
  assign w854[47] = |(datain[123:120] ^ 15);
  assign w854[48] = |(datain[119:116] ^ 14);
  assign w854[49] = |(datain[115:112] ^ 8);
  assign w854[50] = |(datain[111:108] ^ 0);
  assign w854[51] = |(datain[107:104] ^ 0);
  assign w854[52] = |(datain[103:100] ^ 0);
  assign w854[53] = |(datain[99:96] ^ 0);
  assign w854[54] = |(datain[95:92] ^ 5);
  assign w854[55] = |(datain[91:88] ^ 11);
  assign w854[56] = |(datain[87:84] ^ 8);
  assign w854[57] = |(datain[83:80] ^ 9);
  assign w854[58] = |(datain[79:76] ^ 13);
  assign w854[59] = |(datain[75:72] ^ 14);
  assign w854[60] = |(datain[71:68] ^ 8);
  assign w854[61] = |(datain[67:64] ^ 3);
  assign w854[62] = |(datain[63:60] ^ 12);
  assign w854[63] = |(datain[59:56] ^ 3);
  assign w854[64] = |(datain[55:52] ^ 1);
  assign w854[65] = |(datain[51:48] ^ 14);
  assign w854[66] = |(datain[47:44] ^ 8);
  assign w854[67] = |(datain[43:40] ^ 11);
  assign w854[68] = |(datain[39:36] ^ 0);
  assign w854[69] = |(datain[35:32] ^ 7);
  assign w854[70] = |(datain[31:28] ^ 12);
  assign w854[71] = |(datain[27:24] ^ 13);
  assign w854[72] = |(datain[23:20] ^ 2);
  assign w854[73] = |(datain[19:16] ^ 1);
  assign w854[74] = |(datain[15:12] ^ 5);
  assign w854[75] = |(datain[11:8] ^ 14);
  assign comp[854] = ~(|w854);
  wire [76-1:0] w855;
  assign w855[0] = |(datain[311:308] ^ 11);
  assign w855[1] = |(datain[307:304] ^ 9);
  assign w855[2] = |(datain[303:300] ^ 0);
  assign w855[3] = |(datain[299:296] ^ 1);
  assign w855[4] = |(datain[295:292] ^ 0);
  assign w855[5] = |(datain[291:288] ^ 0);
  assign w855[6] = |(datain[287:284] ^ 11);
  assign w855[7] = |(datain[283:280] ^ 11);
  assign w855[8] = |(datain[279:276] ^ 0);
  assign w855[9] = |(datain[275:272] ^ 0);
  assign w855[10] = |(datain[271:268] ^ 0);
  assign w855[11] = |(datain[267:264] ^ 9);
  assign w855[12] = |(datain[263:260] ^ 11);
  assign w855[13] = |(datain[259:256] ^ 8);
  assign w855[14] = |(datain[255:252] ^ 0);
  assign w855[15] = |(datain[251:248] ^ 1);
  assign w855[16] = |(datain[247:244] ^ 0);
  assign w855[17] = |(datain[243:240] ^ 2);
  assign w855[18] = |(datain[239:236] ^ 0);
  assign w855[19] = |(datain[235:232] ^ 14);
  assign w855[20] = |(datain[231:228] ^ 0);
  assign w855[21] = |(datain[227:224] ^ 14);
  assign w855[22] = |(datain[223:220] ^ 0);
  assign w855[23] = |(datain[219:216] ^ 7);
  assign w855[24] = |(datain[215:212] ^ 1);
  assign w855[25] = |(datain[211:208] ^ 15);
  assign w855[26] = |(datain[207:204] ^ 12);
  assign w855[27] = |(datain[203:200] ^ 13);
  assign w855[28] = |(datain[199:196] ^ 1);
  assign w855[29] = |(datain[195:192] ^ 3);
  assign w855[30] = |(datain[191:188] ^ 5);
  assign w855[31] = |(datain[187:184] ^ 1);
  assign w855[32] = |(datain[183:180] ^ 5);
  assign w855[33] = |(datain[179:176] ^ 2);
  assign w855[34] = |(datain[175:172] ^ 5);
  assign w855[35] = |(datain[171:168] ^ 3);
  assign w855[36] = |(datain[167:164] ^ 11);
  assign w855[37] = |(datain[163:160] ^ 9);
  assign w855[38] = |(datain[159:156] ^ 0);
  assign w855[39] = |(datain[155:152] ^ 0);
  assign w855[40] = |(datain[151:148] ^ 0);
  assign w855[41] = |(datain[147:144] ^ 1);
  assign w855[42] = |(datain[143:140] ^ 8);
  assign w855[43] = |(datain[139:136] ^ 11);
  assign w855[44] = |(datain[135:132] ^ 0);
  assign w855[45] = |(datain[131:128] ^ 7);
  assign w855[46] = |(datain[127:124] ^ 4);
  assign w855[47] = |(datain[123:120] ^ 3);
  assign w855[48] = |(datain[119:116] ^ 4);
  assign w855[49] = |(datain[115:112] ^ 3);
  assign w855[50] = |(datain[111:108] ^ 3);
  assign w855[51] = |(datain[107:104] ^ 1);
  assign w855[52] = |(datain[103:100] ^ 0);
  assign w855[53] = |(datain[99:96] ^ 7);
  assign w855[54] = |(datain[95:92] ^ 14);
  assign w855[55] = |(datain[91:88] ^ 2);
  assign w855[56] = |(datain[87:84] ^ 15);
  assign w855[57] = |(datain[83:80] ^ 9);
  assign w855[58] = |(datain[79:76] ^ 5);
  assign w855[59] = |(datain[75:72] ^ 11);
  assign w855[60] = |(datain[71:68] ^ 5);
  assign w855[61] = |(datain[67:64] ^ 10);
  assign w855[62] = |(datain[63:60] ^ 5);
  assign w855[63] = |(datain[59:56] ^ 9);
  assign w855[64] = |(datain[55:52] ^ 11);
  assign w855[65] = |(datain[51:48] ^ 8);
  assign w855[66] = |(datain[47:44] ^ 0);
  assign w855[67] = |(datain[43:40] ^ 1);
  assign w855[68] = |(datain[39:36] ^ 0);
  assign w855[69] = |(datain[35:32] ^ 3);
  assign w855[70] = |(datain[31:28] ^ 12);
  assign w855[71] = |(datain[27:24] ^ 13);
  assign w855[72] = |(datain[23:20] ^ 1);
  assign w855[73] = |(datain[19:16] ^ 3);
  assign w855[74] = |(datain[15:12] ^ 12);
  assign w855[75] = |(datain[11:8] ^ 3);
  assign comp[855] = ~(|w855);
  wire [72-1:0] w856;
  assign w856[0] = |(datain[311:308] ^ 15);
  assign w856[1] = |(datain[307:304] ^ 3);
  assign w856[2] = |(datain[303:300] ^ 10);
  assign w856[3] = |(datain[299:296] ^ 4);
  assign w856[4] = |(datain[295:292] ^ 3);
  assign w856[5] = |(datain[291:288] ^ 14);
  assign w856[6] = |(datain[287:284] ^ 8);
  assign w856[7] = |(datain[283:280] ^ 0);
  assign w856[8] = |(datain[279:276] ^ 8);
  assign w856[9] = |(datain[275:272] ^ 6);
  assign w856[10] = |(datain[271:268] ^ 8);
  assign w856[11] = |(datain[267:264] ^ 10);
  assign w856[12] = |(datain[263:260] ^ 0);
  assign w856[13] = |(datain[259:256] ^ 3);
  assign w856[14] = |(datain[255:252] ^ 0);
  assign w856[15] = |(datain[251:248] ^ 1);
  assign w856[16] = |(datain[247:244] ^ 5);
  assign w856[17] = |(datain[243:240] ^ 11);
  assign w856[18] = |(datain[239:236] ^ 5);
  assign w856[19] = |(datain[235:232] ^ 3);
  assign w856[20] = |(datain[231:228] ^ 11);
  assign w856[21] = |(datain[227:224] ^ 4);
  assign w856[22] = |(datain[223:220] ^ 4);
  assign w856[23] = |(datain[219:216] ^ 0);
  assign w856[24] = |(datain[215:212] ^ 11);
  assign w856[25] = |(datain[211:208] ^ 9);
  assign w856[26] = |(datain[207:204] ^ 0);
  assign w856[27] = |(datain[203:200] ^ 2);
  assign w856[28] = |(datain[199:196] ^ 0);
  assign w856[29] = |(datain[195:192] ^ 0);
  assign w856[30] = |(datain[191:188] ^ 8);
  assign w856[31] = |(datain[187:184] ^ 13);
  assign w856[32] = |(datain[183:180] ^ 9);
  assign w856[33] = |(datain[179:176] ^ 6);
  assign w856[34] = |(datain[175:172] ^ 8);
  assign w856[35] = |(datain[171:168] ^ 10);
  assign w856[36] = |(datain[167:164] ^ 0);
  assign w856[37] = |(datain[163:160] ^ 3);
  assign w856[38] = |(datain[159:156] ^ 12);
  assign w856[39] = |(datain[155:152] ^ 13);
  assign w856[40] = |(datain[151:148] ^ 2);
  assign w856[41] = |(datain[147:144] ^ 1);
  assign w856[42] = |(datain[143:140] ^ 5);
  assign w856[43] = |(datain[139:136] ^ 11);
  assign w856[44] = |(datain[135:132] ^ 5);
  assign w856[45] = |(datain[131:128] ^ 3);
  assign w856[46] = |(datain[127:124] ^ 11);
  assign w856[47] = |(datain[123:120] ^ 4);
  assign w856[48] = |(datain[119:116] ^ 4);
  assign w856[49] = |(datain[115:112] ^ 0);
  assign w856[50] = |(datain[111:108] ^ 11);
  assign w856[51] = |(datain[107:104] ^ 9);
  assign w856[52] = |(datain[103:100] ^ 0);
  assign w856[53] = |(datain[99:96] ^ 4);
  assign w856[54] = |(datain[95:92] ^ 0);
  assign w856[55] = |(datain[91:88] ^ 0);
  assign w856[56] = |(datain[87:84] ^ 8);
  assign w856[57] = |(datain[83:80] ^ 13);
  assign w856[58] = |(datain[79:76] ^ 9);
  assign w856[59] = |(datain[75:72] ^ 6);
  assign w856[60] = |(datain[71:68] ^ 9);
  assign w856[61] = |(datain[67:64] ^ 3);
  assign w856[62] = |(datain[63:60] ^ 0);
  assign w856[63] = |(datain[59:56] ^ 3);
  assign w856[64] = |(datain[55:52] ^ 12);
  assign w856[65] = |(datain[51:48] ^ 13);
  assign w856[66] = |(datain[47:44] ^ 2);
  assign w856[67] = |(datain[43:40] ^ 1);
  assign w856[68] = |(datain[39:36] ^ 5);
  assign w856[69] = |(datain[35:32] ^ 11);
  assign w856[70] = |(datain[31:28] ^ 5);
  assign w856[71] = |(datain[27:24] ^ 3);
  assign comp[856] = ~(|w856);
  wire [74-1:0] w857;
  assign w857[0] = |(datain[311:308] ^ 12);
  assign w857[1] = |(datain[307:304] ^ 9);
  assign w857[2] = |(datain[303:300] ^ 11);
  assign w857[3] = |(datain[299:296] ^ 10);
  assign w857[4] = |(datain[295:292] ^ 11);
  assign w857[5] = |(datain[291:288] ^ 4);
  assign w857[6] = |(datain[287:284] ^ 0);
  assign w857[7] = |(datain[283:280] ^ 1);
  assign w857[8] = |(datain[279:276] ^ 12);
  assign w857[9] = |(datain[275:272] ^ 13);
  assign w857[10] = |(datain[271:268] ^ 2);
  assign w857[11] = |(datain[267:264] ^ 1);
  assign w857[12] = |(datain[263:260] ^ 7);
  assign w857[13] = |(datain[259:256] ^ 2);
  assign w857[14] = |(datain[255:252] ^ 2);
  assign w857[15] = |(datain[251:248] ^ 6);
  assign w857[16] = |(datain[247:244] ^ 11);
  assign w857[17] = |(datain[243:240] ^ 8);
  assign w857[18] = |(datain[239:236] ^ 0);
  assign w857[19] = |(datain[235:232] ^ 1);
  assign w857[20] = |(datain[231:228] ^ 3);
  assign w857[21] = |(datain[227:224] ^ 13);
  assign w857[22] = |(datain[223:220] ^ 11);
  assign w857[23] = |(datain[219:216] ^ 10);
  assign w857[24] = |(datain[215:212] ^ 9);
  assign w857[25] = |(datain[211:208] ^ 14);
  assign w857[26] = |(datain[207:204] ^ 0);
  assign w857[27] = |(datain[203:200] ^ 0);
  assign w857[28] = |(datain[199:196] ^ 12);
  assign w857[29] = |(datain[195:192] ^ 13);
  assign w857[30] = |(datain[191:188] ^ 2);
  assign w857[31] = |(datain[187:184] ^ 1);
  assign w857[32] = |(datain[183:180] ^ 9);
  assign w857[33] = |(datain[179:176] ^ 3);
  assign w857[34] = |(datain[175:172] ^ 11);
  assign w857[35] = |(datain[171:168] ^ 4);
  assign w857[36] = |(datain[167:164] ^ 4);
  assign w857[37] = |(datain[163:160] ^ 0);
  assign w857[38] = |(datain[159:156] ^ 5);
  assign w857[39] = |(datain[155:152] ^ 0);
  assign w857[40] = |(datain[151:148] ^ 11);
  assign w857[41] = |(datain[147:144] ^ 9);
  assign w857[42] = |(datain[143:140] ^ 3);
  assign w857[43] = |(datain[139:136] ^ 1);
  assign w857[44] = |(datain[135:132] ^ 0);
  assign w857[45] = |(datain[131:128] ^ 0);
  assign w857[46] = |(datain[127:124] ^ 11);
  assign w857[47] = |(datain[123:120] ^ 10);
  assign w857[48] = |(datain[119:116] ^ 0);
  assign w857[49] = |(datain[115:112] ^ 0);
  assign w857[50] = |(datain[111:108] ^ 0);
  assign w857[51] = |(datain[107:104] ^ 1);
  assign w857[52] = |(datain[103:100] ^ 12);
  assign w857[53] = |(datain[99:96] ^ 13);
  assign w857[54] = |(datain[95:92] ^ 2);
  assign w857[55] = |(datain[91:88] ^ 1);
  assign w857[56] = |(datain[87:84] ^ 5);
  assign w857[57] = |(datain[83:80] ^ 8);
  assign w857[58] = |(datain[79:76] ^ 11);
  assign w857[59] = |(datain[75:72] ^ 9);
  assign w857[60] = |(datain[71:68] ^ 8);
  assign w857[61] = |(datain[67:64] ^ 8);
  assign w857[62] = |(datain[63:60] ^ 0);
  assign w857[63] = |(datain[59:56] ^ 0);
  assign w857[64] = |(datain[55:52] ^ 11);
  assign w857[65] = |(datain[51:48] ^ 10);
  assign w857[66] = |(datain[47:44] ^ 12);
  assign w857[67] = |(datain[43:40] ^ 3);
  assign w857[68] = |(datain[39:36] ^ 0);
  assign w857[69] = |(datain[35:32] ^ 1);
  assign w857[70] = |(datain[31:28] ^ 12);
  assign w857[71] = |(datain[27:24] ^ 13);
  assign w857[72] = |(datain[23:20] ^ 2);
  assign w857[73] = |(datain[19:16] ^ 1);
  assign comp[857] = ~(|w857);
  wire [74-1:0] w858;
  assign w858[0] = |(datain[311:308] ^ 11);
  assign w858[1] = |(datain[307:304] ^ 9);
  assign w858[2] = |(datain[303:300] ^ 1);
  assign w858[3] = |(datain[299:296] ^ 9);
  assign w858[4] = |(datain[295:292] ^ 0);
  assign w858[5] = |(datain[291:288] ^ 0);
  assign w858[6] = |(datain[287:284] ^ 10);
  assign w858[7] = |(datain[283:280] ^ 4);
  assign w858[8] = |(datain[279:276] ^ 14);
  assign w858[9] = |(datain[275:272] ^ 2);
  assign w858[10] = |(datain[271:268] ^ 15);
  assign w858[11] = |(datain[267:264] ^ 13);
  assign w858[12] = |(datain[263:260] ^ 11);
  assign w858[13] = |(datain[259:256] ^ 10);
  assign w858[14] = |(datain[255:252] ^ 15);
  assign w858[15] = |(datain[251:248] ^ 2);
  assign w858[16] = |(datain[247:244] ^ 0);
  assign w858[17] = |(datain[243:240] ^ 1);
  assign w858[18] = |(datain[239:236] ^ 15);
  assign w858[19] = |(datain[235:232] ^ 15);
  assign w858[20] = |(datain[231:228] ^ 13);
  assign w858[21] = |(datain[227:224] ^ 2);
  assign w858[22] = |(datain[223:220] ^ 12);
  assign w858[23] = |(datain[219:216] ^ 3);
  assign w858[24] = |(datain[215:212] ^ 5);
  assign w858[25] = |(datain[211:208] ^ 3);
  assign w858[26] = |(datain[207:204] ^ 11);
  assign w858[27] = |(datain[203:200] ^ 10);
  assign w858[28] = |(datain[199:196] ^ 13);
  assign w858[29] = |(datain[195:192] ^ 10);
  assign w858[30] = |(datain[191:188] ^ 0);
  assign w858[31] = |(datain[187:184] ^ 1);
  assign w858[32] = |(datain[183:180] ^ 15);
  assign w858[33] = |(datain[179:176] ^ 15);
  assign w858[34] = |(datain[175:172] ^ 13);
  assign w858[35] = |(datain[171:168] ^ 2);
  assign w858[36] = |(datain[167:164] ^ 5);
  assign w858[37] = |(datain[163:160] ^ 11);
  assign w858[38] = |(datain[159:156] ^ 11);
  assign w858[39] = |(datain[155:152] ^ 4);
  assign w858[40] = |(datain[151:148] ^ 4);
  assign w858[41] = |(datain[147:144] ^ 0);
  assign w858[42] = |(datain[143:140] ^ 11);
  assign w858[43] = |(datain[139:136] ^ 9);
  assign w858[44] = |(datain[135:132] ^ 15);
  assign w858[45] = |(datain[131:128] ^ 2);
  assign w858[46] = |(datain[127:124] ^ 0);
  assign w858[47] = |(datain[123:120] ^ 0);
  assign w858[48] = |(datain[119:116] ^ 11);
  assign w858[49] = |(datain[115:112] ^ 10);
  assign w858[50] = |(datain[111:108] ^ 0);
  assign w858[51] = |(datain[107:104] ^ 0);
  assign w858[52] = |(datain[103:100] ^ 0);
  assign w858[53] = |(datain[99:96] ^ 1);
  assign w858[54] = |(datain[95:92] ^ 12);
  assign w858[55] = |(datain[91:88] ^ 13);
  assign w858[56] = |(datain[87:84] ^ 2);
  assign w858[57] = |(datain[83:80] ^ 1);
  assign w858[58] = |(datain[79:76] ^ 5);
  assign w858[59] = |(datain[75:72] ^ 3);
  assign w858[60] = |(datain[71:68] ^ 11);
  assign w858[61] = |(datain[67:64] ^ 10);
  assign w858[62] = |(datain[63:60] ^ 13);
  assign w858[63] = |(datain[59:56] ^ 10);
  assign w858[64] = |(datain[55:52] ^ 0);
  assign w858[65] = |(datain[51:48] ^ 1);
  assign w858[66] = |(datain[47:44] ^ 15);
  assign w858[67] = |(datain[43:40] ^ 15);
  assign w858[68] = |(datain[39:36] ^ 13);
  assign w858[69] = |(datain[35:32] ^ 2);
  assign w858[70] = |(datain[31:28] ^ 5);
  assign w858[71] = |(datain[27:24] ^ 11);
  assign w858[72] = |(datain[23:20] ^ 12);
  assign w858[73] = |(datain[19:16] ^ 3);
  assign comp[858] = ~(|w858);
  wire [72-1:0] w859;
  assign w859[0] = |(datain[311:308] ^ 11);
  assign w859[1] = |(datain[307:304] ^ 15);
  assign w859[2] = |(datain[303:300] ^ 0);
  assign w859[3] = |(datain[299:296] ^ 0);
  assign w859[4] = |(datain[295:292] ^ 0);
  assign w859[5] = |(datain[291:288] ^ 1);
  assign w859[6] = |(datain[287:284] ^ 10);
  assign w859[7] = |(datain[283:280] ^ 5);
  assign w859[8] = |(datain[279:276] ^ 10);
  assign w859[9] = |(datain[275:272] ^ 5);
  assign w859[10] = |(datain[271:268] ^ 8);
  assign w859[11] = |(datain[267:264] ^ 13);
  assign w859[12] = |(datain[263:260] ^ 9);
  assign w859[13] = |(datain[259:256] ^ 6);
  assign w859[14] = |(datain[255:252] ^ 4);
  assign w859[15] = |(datain[251:248] ^ 1);
  assign w859[16] = |(datain[247:244] ^ 0);
  assign w859[17] = |(datain[243:240] ^ 2);
  assign w859[18] = |(datain[239:236] ^ 11);
  assign w859[19] = |(datain[235:232] ^ 4);
  assign w859[20] = |(datain[231:228] ^ 1);
  assign w859[21] = |(datain[227:224] ^ 10);
  assign w859[22] = |(datain[223:220] ^ 12);
  assign w859[23] = |(datain[219:216] ^ 13);
  assign w859[24] = |(datain[215:212] ^ 2);
  assign w859[25] = |(datain[211:208] ^ 1);
  assign w859[26] = |(datain[207:204] ^ 8);
  assign w859[27] = |(datain[203:200] ^ 13);
  assign w859[28] = |(datain[199:196] ^ 9);
  assign w859[29] = |(datain[195:192] ^ 6);
  assign w859[30] = |(datain[191:188] ^ 15);
  assign w859[31] = |(datain[187:184] ^ 1);
  assign w859[32] = |(datain[183:180] ^ 0);
  assign w859[33] = |(datain[179:176] ^ 1);
  assign w859[34] = |(datain[175:172] ^ 11);
  assign w859[35] = |(datain[171:168] ^ 4);
  assign w859[36] = |(datain[167:164] ^ 4);
  assign w859[37] = |(datain[163:160] ^ 14);
  assign w859[38] = |(datain[159:156] ^ 12);
  assign w859[39] = |(datain[155:152] ^ 13);
  assign w859[40] = |(datain[151:148] ^ 2);
  assign w859[41] = |(datain[147:144] ^ 1);
  assign w859[42] = |(datain[143:140] ^ 7);
  assign w859[43] = |(datain[139:136] ^ 2);
  assign w859[44] = |(datain[135:132] ^ 5);
  assign w859[45] = |(datain[131:128] ^ 14);
  assign w859[46] = |(datain[127:124] ^ 8);
  assign w859[47] = |(datain[123:120] ^ 13);
  assign w859[48] = |(datain[119:116] ^ 9);
  assign w859[49] = |(datain[115:112] ^ 6);
  assign w859[50] = |(datain[111:108] ^ 5);
  assign w859[51] = |(datain[107:104] ^ 15);
  assign w859[52] = |(datain[103:100] ^ 0);
  assign w859[53] = |(datain[99:96] ^ 2);
  assign w859[54] = |(datain[95:92] ^ 11);
  assign w859[55] = |(datain[91:88] ^ 8);
  assign w859[56] = |(datain[87:84] ^ 0);
  assign w859[57] = |(datain[83:80] ^ 2);
  assign w859[58] = |(datain[79:76] ^ 3);
  assign w859[59] = |(datain[75:72] ^ 13);
  assign w859[60] = |(datain[71:68] ^ 12);
  assign w859[61] = |(datain[67:64] ^ 13);
  assign w859[62] = |(datain[63:60] ^ 2);
  assign w859[63] = |(datain[59:56] ^ 1);
  assign w859[64] = |(datain[55:52] ^ 9);
  assign w859[65] = |(datain[51:48] ^ 3);
  assign w859[66] = |(datain[47:44] ^ 11);
  assign w859[67] = |(datain[43:40] ^ 9);
  assign w859[68] = |(datain[39:36] ^ 0);
  assign w859[69] = |(datain[35:32] ^ 4);
  assign w859[70] = |(datain[31:28] ^ 0);
  assign w859[71] = |(datain[27:24] ^ 0);
  assign comp[859] = ~(|w859);
  wire [76-1:0] w860;
  assign w860[0] = |(datain[311:308] ^ 11);
  assign w860[1] = |(datain[307:304] ^ 9);
  assign w860[2] = |(datain[303:300] ^ 14);
  assign w860[3] = |(datain[299:296] ^ 7);
  assign w860[4] = |(datain[295:292] ^ 0);
  assign w860[5] = |(datain[291:288] ^ 3);
  assign w860[6] = |(datain[287:284] ^ 8);
  assign w860[7] = |(datain[283:280] ^ 13);
  assign w860[8] = |(datain[279:276] ^ 9);
  assign w860[9] = |(datain[275:272] ^ 6);
  assign w860[10] = |(datain[271:268] ^ 0);
  assign w860[11] = |(datain[267:264] ^ 10);
  assign w860[12] = |(datain[263:260] ^ 0);
  assign w860[13] = |(datain[259:256] ^ 1);
  assign w860[14] = |(datain[255:252] ^ 12);
  assign w860[15] = |(datain[251:248] ^ 13);
  assign w860[16] = |(datain[247:244] ^ 2);
  assign w860[17] = |(datain[243:240] ^ 1);
  assign w860[18] = |(datain[239:236] ^ 5);
  assign w860[19] = |(datain[235:232] ^ 11);
  assign w860[20] = |(datain[231:228] ^ 5);
  assign w860[21] = |(datain[227:224] ^ 3);
  assign w860[22] = |(datain[223:220] ^ 11);
  assign w860[23] = |(datain[219:216] ^ 8);
  assign w860[24] = |(datain[215:212] ^ 0);
  assign w860[25] = |(datain[211:208] ^ 1);
  assign w860[26] = |(datain[207:204] ^ 5);
  assign w860[27] = |(datain[203:200] ^ 7);
  assign w860[28] = |(datain[199:196] ^ 3);
  assign w860[29] = |(datain[195:192] ^ 14);
  assign w860[30] = |(datain[191:188] ^ 8);
  assign w860[31] = |(datain[187:184] ^ 11);
  assign w860[32] = |(datain[183:180] ^ 8);
  assign w860[33] = |(datain[179:176] ^ 14);
  assign w860[34] = |(datain[175:172] ^ 0);
  assign w860[35] = |(datain[171:168] ^ 4);
  assign w860[36] = |(datain[167:164] ^ 0);
  assign w860[37] = |(datain[163:160] ^ 3);
  assign w860[38] = |(datain[159:156] ^ 3);
  assign w860[39] = |(datain[155:152] ^ 14);
  assign w860[40] = |(datain[151:148] ^ 8);
  assign w860[41] = |(datain[147:144] ^ 11);
  assign w860[42] = |(datain[143:140] ^ 9);
  assign w860[43] = |(datain[139:136] ^ 6);
  assign w860[44] = |(datain[135:132] ^ 0);
  assign w860[45] = |(datain[131:128] ^ 6);
  assign w860[46] = |(datain[127:124] ^ 0);
  assign w860[47] = |(datain[123:120] ^ 3);
  assign w860[48] = |(datain[119:116] ^ 12);
  assign w860[49] = |(datain[115:112] ^ 13);
  assign w860[50] = |(datain[111:108] ^ 2);
  assign w860[51] = |(datain[107:104] ^ 1);
  assign w860[52] = |(datain[103:100] ^ 5);
  assign w860[53] = |(datain[99:96] ^ 11);
  assign w860[54] = |(datain[95:92] ^ 11);
  assign w860[55] = |(datain[91:88] ^ 4);
  assign w860[56] = |(datain[87:84] ^ 3);
  assign w860[57] = |(datain[83:80] ^ 14);
  assign w860[58] = |(datain[79:76] ^ 12);
  assign w860[59] = |(datain[75:72] ^ 13);
  assign w860[60] = |(datain[71:68] ^ 2);
  assign w860[61] = |(datain[67:64] ^ 1);
  assign w860[62] = |(datain[63:60] ^ 6);
  assign w860[63] = |(datain[59:56] ^ 8);
  assign w860[64] = |(datain[55:52] ^ 0);
  assign w860[65] = |(datain[51:48] ^ 1);
  assign w860[66] = |(datain[47:44] ^ 4);
  assign w860[67] = |(datain[43:40] ^ 3);
  assign w860[68] = |(datain[39:36] ^ 5);
  assign w860[69] = |(datain[35:32] ^ 8);
  assign w860[70] = |(datain[31:28] ^ 11);
  assign w860[71] = |(datain[27:24] ^ 10);
  assign w860[72] = |(datain[23:20] ^ 9);
  assign w860[73] = |(datain[19:16] ^ 14);
  assign w860[74] = |(datain[15:12] ^ 0);
  assign w860[75] = |(datain[11:8] ^ 0);
  assign comp[860] = ~(|w860);
  wire [72-1:0] w861;
  assign w861[0] = |(datain[311:308] ^ 14);
  assign w861[1] = |(datain[307:304] ^ 8);
  assign w861[2] = |(datain[303:300] ^ 0);
  assign w861[3] = |(datain[299:296] ^ 0);
  assign w861[4] = |(datain[295:292] ^ 0);
  assign w861[5] = |(datain[291:288] ^ 0);
  assign w861[6] = |(datain[287:284] ^ 12);
  assign w861[7] = |(datain[283:280] ^ 12);
  assign w861[8] = |(datain[279:276] ^ 8);
  assign w861[9] = |(datain[275:272] ^ 11);
  assign w861[10] = |(datain[271:268] ^ 15);
  assign w861[11] = |(datain[267:264] ^ 12);
  assign w861[12] = |(datain[263:260] ^ 3);
  assign w861[13] = |(datain[259:256] ^ 6);
  assign w861[14] = |(datain[255:252] ^ 8);
  assign w861[15] = |(datain[251:248] ^ 11);
  assign w861[16] = |(datain[247:244] ^ 2);
  assign w861[17] = |(datain[243:240] ^ 13);
  assign w861[18] = |(datain[239:236] ^ 8);
  assign w861[19] = |(datain[235:232] ^ 1);
  assign w861[20] = |(datain[231:228] ^ 14);
  assign w861[21] = |(datain[227:224] ^ 13);
  assign w861[22] = |(datain[223:220] ^ 1);
  assign w861[23] = |(datain[219:216] ^ 1);
  assign w861[24] = |(datain[215:212] ^ 0);
  assign w861[25] = |(datain[211:208] ^ 1);
  assign w861[26] = |(datain[207:204] ^ 8);
  assign w861[27] = |(datain[203:200] ^ 3);
  assign w861[28] = |(datain[199:196] ^ 12);
  assign w861[29] = |(datain[195:192] ^ 4);
  assign w861[30] = |(datain[191:188] ^ 0);
  assign w861[31] = |(datain[187:184] ^ 2);
  assign w861[32] = |(datain[183:180] ^ 6);
  assign w861[33] = |(datain[179:176] ^ 0);
  assign w861[34] = |(datain[175:172] ^ 11);
  assign w861[35] = |(datain[171:168] ^ 4);
  assign w861[36] = |(datain[167:164] ^ 2);
  assign w861[37] = |(datain[163:160] ^ 10);
  assign w861[38] = |(datain[159:156] ^ 12);
  assign w861[39] = |(datain[155:152] ^ 13);
  assign w861[40] = |(datain[151:148] ^ 2);
  assign w861[41] = |(datain[147:144] ^ 1);
  assign w861[42] = |(datain[143:140] ^ 8);
  assign w861[43] = |(datain[139:136] ^ 0);
  assign w861[44] = |(datain[135:132] ^ 15);
  assign w861[45] = |(datain[131:128] ^ 10);
  assign w861[46] = |(datain[127:124] ^ 1);
  assign w861[47] = |(datain[123:120] ^ 2);
  assign w861[48] = |(datain[119:116] ^ 7);
  assign w861[49] = |(datain[115:112] ^ 5);
  assign w861[50] = |(datain[111:108] ^ 0);
  assign w861[51] = |(datain[107:104] ^ 7);
  assign w861[52] = |(datain[103:100] ^ 11);
  assign w861[53] = |(datain[99:96] ^ 9);
  assign w861[54] = |(datain[95:92] ^ 15);
  assign w861[55] = |(datain[91:88] ^ 15);
  assign w861[56] = |(datain[87:84] ^ 15);
  assign w861[57] = |(datain[83:80] ^ 15);
  assign w861[58] = |(datain[79:76] ^ 11);
  assign w861[59] = |(datain[75:72] ^ 0);
  assign w861[60] = |(datain[71:68] ^ 0);
  assign w861[61] = |(datain[67:64] ^ 2);
  assign w861[62] = |(datain[63:60] ^ 12);
  assign w861[63] = |(datain[59:56] ^ 13);
  assign w861[64] = |(datain[55:52] ^ 2);
  assign w861[65] = |(datain[51:48] ^ 6);
  assign w861[66] = |(datain[47:44] ^ 6);
  assign w861[67] = |(datain[43:40] ^ 1);
  assign w861[68] = |(datain[39:36] ^ 14);
  assign w861[69] = |(datain[35:32] ^ 8);
  assign w861[70] = |(datain[31:28] ^ 0);
  assign w861[71] = |(datain[27:24] ^ 5);
  assign comp[861] = ~(|w861);
  wire [74-1:0] w862;
  assign w862[0] = |(datain[311:308] ^ 11);
  assign w862[1] = |(datain[307:304] ^ 4);
  assign w862[2] = |(datain[303:300] ^ 4);
  assign w862[3] = |(datain[299:296] ^ 0);
  assign w862[4] = |(datain[295:292] ^ 11);
  assign w862[5] = |(datain[291:288] ^ 9);
  assign w862[6] = |(datain[287:284] ^ 14);
  assign w862[7] = |(datain[283:280] ^ 7);
  assign w862[8] = |(datain[279:276] ^ 0);
  assign w862[9] = |(datain[275:272] ^ 3);
  assign w862[10] = |(datain[271:268] ^ 8);
  assign w862[11] = |(datain[267:264] ^ 13);
  assign w862[12] = |(datain[263:260] ^ 9);
  assign w862[13] = |(datain[259:256] ^ 6);
  assign w862[14] = |(datain[255:252] ^ 0);
  assign w862[15] = |(datain[251:248] ^ 9);
  assign w862[16] = |(datain[247:244] ^ 0);
  assign w862[17] = |(datain[243:240] ^ 1);
  assign w862[18] = |(datain[239:236] ^ 12);
  assign w862[19] = |(datain[235:232] ^ 13);
  assign w862[20] = |(datain[231:228] ^ 2);
  assign w862[21] = |(datain[227:224] ^ 1);
  assign w862[22] = |(datain[223:220] ^ 5);
  assign w862[23] = |(datain[219:216] ^ 11);
  assign w862[24] = |(datain[215:212] ^ 5);
  assign w862[25] = |(datain[211:208] ^ 3);
  assign w862[26] = |(datain[207:204] ^ 11);
  assign w862[27] = |(datain[203:200] ^ 8);
  assign w862[28] = |(datain[199:196] ^ 0);
  assign w862[29] = |(datain[195:192] ^ 1);
  assign w862[30] = |(datain[191:188] ^ 5);
  assign w862[31] = |(datain[187:184] ^ 7);
  assign w862[32] = |(datain[183:180] ^ 3);
  assign w862[33] = |(datain[179:176] ^ 14);
  assign w862[34] = |(datain[175:172] ^ 8);
  assign w862[35] = |(datain[171:168] ^ 11);
  assign w862[36] = |(datain[167:164] ^ 8);
  assign w862[37] = |(datain[163:160] ^ 14);
  assign w862[38] = |(datain[159:156] ^ 4);
  assign w862[39] = |(datain[155:152] ^ 0);
  assign w862[40] = |(datain[151:148] ^ 0);
  assign w862[41] = |(datain[147:144] ^ 3);
  assign w862[42] = |(datain[143:140] ^ 3);
  assign w862[43] = |(datain[139:136] ^ 14);
  assign w862[44] = |(datain[135:132] ^ 8);
  assign w862[45] = |(datain[131:128] ^ 11);
  assign w862[46] = |(datain[127:124] ^ 9);
  assign w862[47] = |(datain[123:120] ^ 6);
  assign w862[48] = |(datain[119:116] ^ 4);
  assign w862[49] = |(datain[115:112] ^ 2);
  assign w862[50] = |(datain[111:108] ^ 0);
  assign w862[51] = |(datain[107:104] ^ 3);
  assign w862[52] = |(datain[103:100] ^ 12);
  assign w862[53] = |(datain[99:96] ^ 13);
  assign w862[54] = |(datain[95:92] ^ 2);
  assign w862[55] = |(datain[91:88] ^ 1);
  assign w862[56] = |(datain[87:84] ^ 5);
  assign w862[57] = |(datain[83:80] ^ 11);
  assign w862[58] = |(datain[79:76] ^ 11);
  assign w862[59] = |(datain[75:72] ^ 4);
  assign w862[60] = |(datain[71:68] ^ 3);
  assign w862[61] = |(datain[67:64] ^ 14);
  assign w862[62] = |(datain[63:60] ^ 12);
  assign w862[63] = |(datain[59:56] ^ 13);
  assign w862[64] = |(datain[55:52] ^ 2);
  assign w862[65] = |(datain[51:48] ^ 1);
  assign w862[66] = |(datain[47:44] ^ 6);
  assign w862[67] = |(datain[43:40] ^ 8);
  assign w862[68] = |(datain[39:36] ^ 0);
  assign w862[69] = |(datain[35:32] ^ 1);
  assign w862[70] = |(datain[31:28] ^ 4);
  assign w862[71] = |(datain[27:24] ^ 3);
  assign w862[72] = |(datain[23:20] ^ 5);
  assign w862[73] = |(datain[19:16] ^ 8);
  assign comp[862] = ~(|w862);
  wire [76-1:0] w863;
  assign w863[0] = |(datain[311:308] ^ 5);
  assign w863[1] = |(datain[307:304] ^ 11);
  assign w863[2] = |(datain[303:300] ^ 5);
  assign w863[3] = |(datain[299:296] ^ 3);
  assign w863[4] = |(datain[295:292] ^ 14);
  assign w863[5] = |(datain[291:288] ^ 8);
  assign w863[6] = |(datain[287:284] ^ 6);
  assign w863[7] = |(datain[283:280] ^ 8);
  assign w863[8] = |(datain[279:276] ^ 15);
  assign w863[9] = |(datain[275:272] ^ 14);
  assign w863[10] = |(datain[271:268] ^ 11);
  assign w863[11] = |(datain[267:264] ^ 4);
  assign w863[12] = |(datain[263:260] ^ 4);
  assign w863[13] = |(datain[259:256] ^ 0);
  assign w863[14] = |(datain[255:252] ^ 11);
  assign w863[15] = |(datain[251:248] ^ 9);
  assign w863[16] = |(datain[247:244] ^ 14);
  assign w863[17] = |(datain[243:240] ^ 7);
  assign w863[18] = |(datain[239:236] ^ 0);
  assign w863[19] = |(datain[235:232] ^ 3);
  assign w863[20] = |(datain[231:228] ^ 8);
  assign w863[21] = |(datain[227:224] ^ 13);
  assign w863[22] = |(datain[223:220] ^ 9);
  assign w863[23] = |(datain[219:216] ^ 6);
  assign w863[24] = |(datain[215:212] ^ 0);
  assign w863[25] = |(datain[211:208] ^ 10);
  assign w863[26] = |(datain[207:204] ^ 0);
  assign w863[27] = |(datain[203:200] ^ 1);
  assign w863[28] = |(datain[199:196] ^ 12);
  assign w863[29] = |(datain[195:192] ^ 13);
  assign w863[30] = |(datain[191:188] ^ 2);
  assign w863[31] = |(datain[187:184] ^ 1);
  assign w863[32] = |(datain[183:180] ^ 5);
  assign w863[33] = |(datain[179:176] ^ 11);
  assign w863[34] = |(datain[175:172] ^ 5);
  assign w863[35] = |(datain[171:168] ^ 3);
  assign w863[36] = |(datain[167:164] ^ 11);
  assign w863[37] = |(datain[163:160] ^ 8);
  assign w863[38] = |(datain[159:156] ^ 0);
  assign w863[39] = |(datain[155:152] ^ 1);
  assign w863[40] = |(datain[151:148] ^ 5);
  assign w863[41] = |(datain[147:144] ^ 7);
  assign w863[42] = |(datain[143:140] ^ 3);
  assign w863[43] = |(datain[139:136] ^ 14);
  assign w863[44] = |(datain[135:132] ^ 8);
  assign w863[45] = |(datain[131:128] ^ 11);
  assign w863[46] = |(datain[127:124] ^ 8);
  assign w863[47] = |(datain[123:120] ^ 14);
  assign w863[48] = |(datain[119:116] ^ 9);
  assign w863[49] = |(datain[115:112] ^ 8);
  assign w863[50] = |(datain[111:108] ^ 0);
  assign w863[51] = |(datain[107:104] ^ 3);
  assign w863[52] = |(datain[103:100] ^ 3);
  assign w863[53] = |(datain[99:96] ^ 14);
  assign w863[54] = |(datain[95:92] ^ 8);
  assign w863[55] = |(datain[91:88] ^ 11);
  assign w863[56] = |(datain[87:84] ^ 9);
  assign w863[57] = |(datain[83:80] ^ 6);
  assign w863[58] = |(datain[79:76] ^ 9);
  assign w863[59] = |(datain[75:72] ^ 10);
  assign w863[60] = |(datain[71:68] ^ 0);
  assign w863[61] = |(datain[67:64] ^ 3);
  assign w863[62] = |(datain[63:60] ^ 12);
  assign w863[63] = |(datain[59:56] ^ 13);
  assign w863[64] = |(datain[55:52] ^ 2);
  assign w863[65] = |(datain[51:48] ^ 1);
  assign w863[66] = |(datain[47:44] ^ 5);
  assign w863[67] = |(datain[43:40] ^ 11);
  assign w863[68] = |(datain[39:36] ^ 11);
  assign w863[69] = |(datain[35:32] ^ 4);
  assign w863[70] = |(datain[31:28] ^ 3);
  assign w863[71] = |(datain[27:24] ^ 14);
  assign w863[72] = |(datain[23:20] ^ 12);
  assign w863[73] = |(datain[19:16] ^ 13);
  assign w863[74] = |(datain[15:12] ^ 2);
  assign w863[75] = |(datain[11:8] ^ 1);
  assign comp[863] = ~(|w863);
  wire [76-1:0] w864;
  assign w864[0] = |(datain[311:308] ^ 5);
  assign w864[1] = |(datain[307:304] ^ 11);
  assign w864[2] = |(datain[303:300] ^ 5);
  assign w864[3] = |(datain[299:296] ^ 3);
  assign w864[4] = |(datain[295:292] ^ 14);
  assign w864[5] = |(datain[291:288] ^ 8);
  assign w864[6] = |(datain[287:284] ^ 6);
  assign w864[7] = |(datain[283:280] ^ 9);
  assign w864[8] = |(datain[279:276] ^ 15);
  assign w864[9] = |(datain[275:272] ^ 14);
  assign w864[10] = |(datain[271:268] ^ 11);
  assign w864[11] = |(datain[267:264] ^ 4);
  assign w864[12] = |(datain[263:260] ^ 4);
  assign w864[13] = |(datain[259:256] ^ 0);
  assign w864[14] = |(datain[255:252] ^ 11);
  assign w864[15] = |(datain[251:248] ^ 9);
  assign w864[16] = |(datain[247:244] ^ 14);
  assign w864[17] = |(datain[243:240] ^ 7);
  assign w864[18] = |(datain[239:236] ^ 0);
  assign w864[19] = |(datain[235:232] ^ 3);
  assign w864[20] = |(datain[231:228] ^ 8);
  assign w864[21] = |(datain[227:224] ^ 13);
  assign w864[22] = |(datain[223:220] ^ 9);
  assign w864[23] = |(datain[219:216] ^ 6);
  assign w864[24] = |(datain[215:212] ^ 0);
  assign w864[25] = |(datain[211:208] ^ 9);
  assign w864[26] = |(datain[207:204] ^ 0);
  assign w864[27] = |(datain[203:200] ^ 1);
  assign w864[28] = |(datain[199:196] ^ 12);
  assign w864[29] = |(datain[195:192] ^ 13);
  assign w864[30] = |(datain[191:188] ^ 2);
  assign w864[31] = |(datain[187:184] ^ 1);
  assign w864[32] = |(datain[183:180] ^ 5);
  assign w864[33] = |(datain[179:176] ^ 11);
  assign w864[34] = |(datain[175:172] ^ 5);
  assign w864[35] = |(datain[171:168] ^ 3);
  assign w864[36] = |(datain[167:164] ^ 11);
  assign w864[37] = |(datain[163:160] ^ 8);
  assign w864[38] = |(datain[159:156] ^ 0);
  assign w864[39] = |(datain[155:152] ^ 1);
  assign w864[40] = |(datain[151:148] ^ 5);
  assign w864[41] = |(datain[147:144] ^ 7);
  assign w864[42] = |(datain[143:140] ^ 3);
  assign w864[43] = |(datain[139:136] ^ 14);
  assign w864[44] = |(datain[135:132] ^ 8);
  assign w864[45] = |(datain[131:128] ^ 11);
  assign w864[46] = |(datain[127:124] ^ 8);
  assign w864[47] = |(datain[123:120] ^ 14);
  assign w864[48] = |(datain[119:116] ^ 11);
  assign w864[49] = |(datain[115:112] ^ 7);
  assign w864[50] = |(datain[111:108] ^ 0);
  assign w864[51] = |(datain[107:104] ^ 3);
  assign w864[52] = |(datain[103:100] ^ 3);
  assign w864[53] = |(datain[99:96] ^ 14);
  assign w864[54] = |(datain[95:92] ^ 8);
  assign w864[55] = |(datain[91:88] ^ 11);
  assign w864[56] = |(datain[87:84] ^ 9);
  assign w864[57] = |(datain[83:80] ^ 6);
  assign w864[58] = |(datain[79:76] ^ 11);
  assign w864[59] = |(datain[75:72] ^ 9);
  assign w864[60] = |(datain[71:68] ^ 0);
  assign w864[61] = |(datain[67:64] ^ 3);
  assign w864[62] = |(datain[63:60] ^ 12);
  assign w864[63] = |(datain[59:56] ^ 13);
  assign w864[64] = |(datain[55:52] ^ 2);
  assign w864[65] = |(datain[51:48] ^ 1);
  assign w864[66] = |(datain[47:44] ^ 5);
  assign w864[67] = |(datain[43:40] ^ 11);
  assign w864[68] = |(datain[39:36] ^ 11);
  assign w864[69] = |(datain[35:32] ^ 4);
  assign w864[70] = |(datain[31:28] ^ 3);
  assign w864[71] = |(datain[27:24] ^ 14);
  assign w864[72] = |(datain[23:20] ^ 12);
  assign w864[73] = |(datain[19:16] ^ 13);
  assign w864[74] = |(datain[15:12] ^ 2);
  assign w864[75] = |(datain[11:8] ^ 1);
  assign comp[864] = ~(|w864);
  wire [74-1:0] w865;
  assign w865[0] = |(datain[311:308] ^ 11);
  assign w865[1] = |(datain[307:304] ^ 10);
  assign w865[2] = |(datain[303:300] ^ 8);
  assign w865[3] = |(datain[299:296] ^ 0);
  assign w865[4] = |(datain[295:292] ^ 0);
  assign w865[5] = |(datain[291:288] ^ 0);
  assign w865[6] = |(datain[287:284] ^ 11);
  assign w865[7] = |(datain[283:280] ^ 9);
  assign w865[8] = |(datain[279:276] ^ 0);
  assign w865[9] = |(datain[275:272] ^ 1);
  assign w865[10] = |(datain[271:268] ^ 0);
  assign w865[11] = |(datain[267:264] ^ 0);
  assign w865[12] = |(datain[263:260] ^ 11);
  assign w865[13] = |(datain[259:256] ^ 11);
  assign w865[14] = |(datain[255:252] ^ 0);
  assign w865[15] = |(datain[251:248] ^ 2);
  assign w865[16] = |(datain[247:244] ^ 0);
  assign w865[17] = |(datain[243:240] ^ 1);
  assign w865[18] = |(datain[239:236] ^ 12);
  assign w865[19] = |(datain[235:232] ^ 7);
  assign w865[20] = |(datain[231:228] ^ 4);
  assign w865[21] = |(datain[227:224] ^ 7);
  assign w865[22] = |(datain[223:220] ^ 1);
  assign w865[23] = |(datain[219:216] ^ 10);
  assign w865[24] = |(datain[215:212] ^ 0);
  assign w865[25] = |(datain[211:208] ^ 0);
  assign w865[26] = |(datain[207:204] ^ 0);
  assign w865[27] = |(datain[203:200] ^ 0);
  assign w865[28] = |(datain[199:196] ^ 12);
  assign w865[29] = |(datain[195:192] ^ 13);
  assign w865[30] = |(datain[191:188] ^ 1);
  assign w865[31] = |(datain[187:184] ^ 3);
  assign w865[32] = |(datain[183:180] ^ 14);
  assign w865[33] = |(datain[179:176] ^ 11);
  assign w865[34] = |(datain[175:172] ^ 1);
  assign w865[35] = |(datain[171:168] ^ 10);
  assign w865[36] = |(datain[167:164] ^ 11);
  assign w865[37] = |(datain[163:160] ^ 4);
  assign w865[38] = |(datain[159:156] ^ 0);
  assign w865[39] = |(datain[155:152] ^ 9);
  assign w865[40] = |(datain[151:148] ^ 11);
  assign w865[41] = |(datain[147:144] ^ 10);
  assign w865[42] = |(datain[143:140] ^ 1);
  assign w865[43] = |(datain[139:136] ^ 4);
  assign w865[44] = |(datain[135:132] ^ 0);
  assign w865[45] = |(datain[131:128] ^ 2);
  assign w865[46] = |(datain[127:124] ^ 8);
  assign w865[47] = |(datain[123:120] ^ 11);
  assign w865[48] = |(datain[119:116] ^ 15);
  assign w865[49] = |(datain[115:112] ^ 2);
  assign w865[50] = |(datain[111:108] ^ 11);
  assign w865[51] = |(datain[107:104] ^ 9);
  assign w865[52] = |(datain[103:100] ^ 2);
  assign w865[53] = |(datain[99:96] ^ 11);
  assign w865[54] = |(datain[95:92] ^ 0);
  assign w865[55] = |(datain[91:88] ^ 0);
  assign w865[56] = |(datain[87:84] ^ 5);
  assign w865[57] = |(datain[83:80] ^ 1);
  assign w865[58] = |(datain[79:76] ^ 15);
  assign w865[59] = |(datain[75:72] ^ 14);
  assign w865[60] = |(datain[71:68] ^ 0);
  assign w865[61] = |(datain[67:64] ^ 12);
  assign w865[62] = |(datain[63:60] ^ 4);
  assign w865[63] = |(datain[59:56] ^ 6);
  assign w865[64] = |(datain[55:52] ^ 14);
  assign w865[65] = |(datain[51:48] ^ 2);
  assign w865[66] = |(datain[47:44] ^ 15);
  assign w865[67] = |(datain[43:40] ^ 11);
  assign w865[68] = |(datain[39:36] ^ 12);
  assign w865[69] = |(datain[35:32] ^ 13);
  assign w865[70] = |(datain[31:28] ^ 2);
  assign w865[71] = |(datain[27:24] ^ 1);
  assign w865[72] = |(datain[23:20] ^ 5);
  assign w865[73] = |(datain[19:16] ^ 9);
  assign comp[865] = ~(|w865);
  wire [74-1:0] w866;
  assign w866[0] = |(datain[311:308] ^ 8);
  assign w866[1] = |(datain[307:304] ^ 1);
  assign w866[2] = |(datain[303:300] ^ 14);
  assign w866[3] = |(datain[299:296] ^ 14);
  assign w866[4] = |(datain[295:292] ^ 5);
  assign w866[5] = |(datain[291:288] ^ 0);
  assign w866[6] = |(datain[287:284] ^ 0);
  assign w866[7] = |(datain[283:280] ^ 1);
  assign w866[8] = |(datain[279:276] ^ 11);
  assign w866[9] = |(datain[275:272] ^ 8);
  assign w866[10] = |(datain[271:268] ^ 12);
  assign w866[11] = |(datain[267:264] ^ 13);
  assign w866[12] = |(datain[263:260] ^ 10);
  assign w866[13] = |(datain[259:256] ^ 11);
  assign w866[14] = |(datain[255:252] ^ 8);
  assign w866[15] = |(datain[251:248] ^ 11);
  assign w866[16] = |(datain[247:244] ^ 0);
  assign w866[17] = |(datain[243:240] ^ 12);
  assign w866[18] = |(datain[239:236] ^ 3);
  assign w866[19] = |(datain[235:232] ^ 1);
  assign w866[20] = |(datain[231:228] ^ 13);
  assign w866[21] = |(datain[227:224] ^ 2);
  assign w866[22] = |(datain[223:220] ^ 3);
  assign w866[23] = |(datain[219:216] ^ 1);
  assign w866[24] = |(datain[215:212] ^ 12);
  assign w866[25] = |(datain[211:208] ^ 1);
  assign w866[26] = |(datain[207:204] ^ 4);
  assign w866[27] = |(datain[203:200] ^ 8);
  assign w866[28] = |(datain[199:196] ^ 0);
  assign w866[29] = |(datain[195:192] ^ 1);
  assign w866[30] = |(datain[191:188] ^ 12);
  assign w866[31] = |(datain[187:184] ^ 0);
  assign w866[32] = |(datain[183:180] ^ 8);
  assign w866[33] = |(datain[179:176] ^ 10);
  assign w866[34] = |(datain[175:172] ^ 15);
  assign w866[35] = |(datain[171:168] ^ 5);
  assign w866[36] = |(datain[167:164] ^ 8);
  assign w866[37] = |(datain[163:160] ^ 10);
  assign w866[38] = |(datain[159:156] ^ 13);
  assign w866[39] = |(datain[155:152] ^ 1);
  assign w866[40] = |(datain[151:148] ^ 8);
  assign w866[41] = |(datain[147:144] ^ 9);
  assign w866[42] = |(datain[143:140] ^ 1);
  assign w866[43] = |(datain[139:136] ^ 4);
  assign w866[44] = |(datain[135:132] ^ 4);
  assign w866[45] = |(datain[131:128] ^ 6);
  assign w866[46] = |(datain[127:124] ^ 8);
  assign w866[47] = |(datain[123:120] ^ 1);
  assign w866[48] = |(datain[119:116] ^ 15);
  assign w866[49] = |(datain[115:112] ^ 14);
  assign w866[50] = |(datain[111:108] ^ 10);
  assign w866[51] = |(datain[107:104] ^ 5);
  assign w866[52] = |(datain[103:100] ^ 1);
  assign w866[53] = |(datain[99:96] ^ 3);
  assign w866[54] = |(datain[95:92] ^ 7);
  assign w866[55] = |(datain[91:88] ^ 5);
  assign w866[56] = |(datain[87:84] ^ 14);
  assign w866[57] = |(datain[83:80] ^ 10);
  assign w866[58] = |(datain[79:76] ^ 8);
  assign w866[59] = |(datain[75:72] ^ 12);
  assign w866[60] = |(datain[71:68] ^ 13);
  assign w866[61] = |(datain[67:64] ^ 9);
  assign w866[62] = |(datain[63:60] ^ 8);
  assign w866[63] = |(datain[59:56] ^ 1);
  assign w866[64] = |(datain[55:52] ^ 12);
  assign w866[65] = |(datain[51:48] ^ 1);
  assign w866[66] = |(datain[47:44] ^ 1);
  assign w866[67] = |(datain[43:40] ^ 0);
  assign w866[68] = |(datain[39:36] ^ 0);
  assign w866[69] = |(datain[35:32] ^ 0);
  assign w866[70] = |(datain[31:28] ^ 8);
  assign w866[71] = |(datain[27:24] ^ 14);
  assign w866[72] = |(datain[23:20] ^ 12);
  assign w866[73] = |(datain[19:16] ^ 1);
  assign comp[866] = ~(|w866);
  wire [42-1:0] w867;
  assign w867[0] = |(datain[311:308] ^ 13);
  assign w867[1] = |(datain[307:304] ^ 8);
  assign w867[2] = |(datain[303:300] ^ 11);
  assign w867[3] = |(datain[299:296] ^ 8);
  assign w867[4] = |(datain[295:292] ^ 0);
  assign w867[5] = |(datain[291:288] ^ 0);
  assign w867[6] = |(datain[287:284] ^ 4);
  assign w867[7] = |(datain[283:280] ^ 0);
  assign w867[8] = |(datain[279:276] ^ 11);
  assign w867[9] = |(datain[275:272] ^ 9);
  assign w867[10] = |(datain[271:268] ^ 11);
  assign w867[11] = |(datain[267:264] ^ 0);
  assign w867[12] = |(datain[263:260] ^ 0);
  assign w867[13] = |(datain[259:256] ^ 1);
  assign w867[14] = |(datain[255:252] ^ 3);
  assign w867[15] = |(datain[251:248] ^ 3);
  assign w867[16] = |(datain[247:244] ^ 13);
  assign w867[17] = |(datain[243:240] ^ 2);
  assign w867[18] = |(datain[239:236] ^ 12);
  assign w867[19] = |(datain[235:232] ^ 13);
  assign w867[20] = |(datain[231:228] ^ 2);
  assign w867[21] = |(datain[227:224] ^ 1);
  assign w867[22] = |(datain[223:220] ^ 7);
  assign w867[23] = |(datain[219:216] ^ 2);
  assign w867[24] = |(datain[215:212] ^ 1);
  assign w867[25] = |(datain[211:208] ^ 11);
  assign w867[26] = |(datain[207:204] ^ 11);
  assign w867[27] = |(datain[203:200] ^ 8);
  assign w867[28] = |(datain[199:196] ^ 0);
  assign w867[29] = |(datain[195:192] ^ 0);
  assign w867[30] = |(datain[191:188] ^ 4);
  assign w867[31] = |(datain[187:184] ^ 2);
  assign w867[32] = |(datain[183:180] ^ 3);
  assign w867[33] = |(datain[179:176] ^ 3);
  assign w867[34] = |(datain[175:172] ^ 12);
  assign w867[35] = |(datain[171:168] ^ 9);
  assign w867[36] = |(datain[167:164] ^ 3);
  assign w867[37] = |(datain[163:160] ^ 3);
  assign w867[38] = |(datain[159:156] ^ 13);
  assign w867[39] = |(datain[155:152] ^ 2);
  assign w867[40] = |(datain[151:148] ^ 12);
  assign w867[41] = |(datain[147:144] ^ 13);
  assign comp[867] = ~(|w867);
  wire [46-1:0] w868;
  assign w868[0] = |(datain[311:308] ^ 14);
  assign w868[1] = |(datain[307:304] ^ 2);
  assign w868[2] = |(datain[303:300] ^ 11);
  assign w868[3] = |(datain[299:296] ^ 15);
  assign w868[4] = |(datain[295:292] ^ 8);
  assign w868[5] = |(datain[291:288] ^ 14);
  assign w868[6] = |(datain[287:284] ^ 12);
  assign w868[7] = |(datain[283:280] ^ 0);
  assign w868[8] = |(datain[279:276] ^ 8);
  assign w868[9] = |(datain[275:272] ^ 9);
  assign w868[10] = |(datain[271:268] ^ 13);
  assign w868[11] = |(datain[267:264] ^ 14);
  assign w868[12] = |(datain[263:260] ^ 3);
  assign w868[13] = |(datain[259:256] ^ 3);
  assign w868[14] = |(datain[255:252] ^ 15);
  assign w868[15] = |(datain[251:248] ^ 15);
  assign w868[16] = |(datain[247:244] ^ 11);
  assign w868[17] = |(datain[243:240] ^ 9);
  assign w868[18] = |(datain[239:236] ^ 13);
  assign w868[19] = |(datain[235:232] ^ 13);
  assign w868[20] = |(datain[231:228] ^ 0);
  assign w868[21] = |(datain[227:224] ^ 1);
  assign w868[22] = |(datain[223:220] ^ 15);
  assign w868[23] = |(datain[219:216] ^ 3);
  assign w868[24] = |(datain[215:212] ^ 10);
  assign w868[25] = |(datain[211:208] ^ 4);
  assign w868[26] = |(datain[207:204] ^ 8);
  assign w868[27] = |(datain[203:200] ^ 9);
  assign w868[28] = |(datain[199:196] ^ 13);
  assign w868[29] = |(datain[195:192] ^ 14);
  assign w868[30] = |(datain[191:188] ^ 3);
  assign w868[31] = |(datain[187:184] ^ 3);
  assign w868[32] = |(datain[183:180] ^ 15);
  assign w868[33] = |(datain[179:176] ^ 15);
  assign w868[34] = |(datain[175:172] ^ 11);
  assign w868[35] = |(datain[171:168] ^ 9);
  assign w868[36] = |(datain[167:164] ^ 13);
  assign w868[37] = |(datain[163:160] ^ 13);
  assign w868[38] = |(datain[159:156] ^ 0);
  assign w868[39] = |(datain[155:152] ^ 1);
  assign w868[40] = |(datain[151:148] ^ 15);
  assign w868[41] = |(datain[147:144] ^ 3);
  assign w868[42] = |(datain[143:140] ^ 10);
  assign w868[43] = |(datain[139:136] ^ 6);
  assign w868[44] = |(datain[135:132] ^ 7);
  assign w868[45] = |(datain[131:128] ^ 4);
  assign comp[868] = ~(|w868);
  wire [56-1:0] w869;
  assign w869[0] = |(datain[311:308] ^ 11);
  assign w869[1] = |(datain[307:304] ^ 12);
  assign w869[2] = |(datain[303:300] ^ 15);
  assign w869[3] = |(datain[299:296] ^ 10);
  assign w869[4] = |(datain[295:292] ^ 11);
  assign w869[5] = |(datain[291:288] ^ 4);
  assign w869[6] = |(datain[287:284] ^ 8);
  assign w869[7] = |(datain[283:280] ^ 13);
  assign w869[8] = |(datain[279:276] ^ 12);
  assign w869[9] = |(datain[275:272] ^ 4);
  assign w869[10] = |(datain[271:268] ^ 12);
  assign w869[11] = |(datain[267:264] ^ 9);
  assign w869[12] = |(datain[263:260] ^ 2);
  assign w869[13] = |(datain[259:256] ^ 11);
  assign w869[14] = |(datain[255:252] ^ 14);
  assign w869[15] = |(datain[251:248] ^ 15);
  assign w869[16] = |(datain[247:244] ^ 0);
  assign w869[17] = |(datain[243:240] ^ 4);
  assign w869[18] = |(datain[239:236] ^ 0);
  assign w869[19] = |(datain[235:232] ^ 10);
  assign w869[20] = |(datain[231:228] ^ 1);
  assign w869[21] = |(datain[227:224] ^ 11);
  assign w869[22] = |(datain[223:220] ^ 12);
  assign w869[23] = |(datain[219:216] ^ 2);
  assign w869[24] = |(datain[215:212] ^ 0);
  assign w869[25] = |(datain[211:208] ^ 2);
  assign w869[26] = |(datain[207:204] ^ 14);
  assign w869[27] = |(datain[203:200] ^ 12);
  assign w869[28] = |(datain[199:196] ^ 0);
  assign w869[29] = |(datain[195:192] ^ 14);
  assign w869[30] = |(datain[191:188] ^ 0);
  assign w869[31] = |(datain[187:184] ^ 4);
  assign w869[32] = |(datain[183:180] ^ 14);
  assign w869[33] = |(datain[179:176] ^ 12);
  assign w869[34] = |(datain[175:172] ^ 13);
  assign w869[35] = |(datain[171:168] ^ 12);
  assign w869[36] = |(datain[167:164] ^ 0);
  assign w869[37] = |(datain[163:160] ^ 4);
  assign w869[38] = |(datain[159:156] ^ 11);
  assign w869[39] = |(datain[155:152] ^ 12);
  assign w869[40] = |(datain[151:148] ^ 0);
  assign w869[41] = |(datain[147:144] ^ 4);
  assign w869[42] = |(datain[143:140] ^ 1);
  assign w869[43] = |(datain[139:136] ^ 6);
  assign w869[44] = |(datain[135:132] ^ 12);
  assign w869[45] = |(datain[131:128] ^ 9);
  assign w869[46] = |(datain[127:124] ^ 2);
  assign w869[47] = |(datain[123:120] ^ 11);
  assign w869[48] = |(datain[119:116] ^ 15);
  assign w869[49] = |(datain[115:112] ^ 10);
  assign w869[50] = |(datain[111:108] ^ 12);
  assign w869[51] = |(datain[107:104] ^ 4);
  assign w869[52] = |(datain[103:100] ^ 7);
  assign w869[53] = |(datain[99:96] ^ 1);
  assign w869[54] = |(datain[95:92] ^ 0);
  assign w869[55] = |(datain[91:88] ^ 12);
  assign comp[869] = ~(|w869);
  wire [64-1:0] w870;
  assign w870[0] = |(datain[311:308] ^ 11);
  assign w870[1] = |(datain[307:304] ^ 0);
  assign w870[2] = |(datain[303:300] ^ 8);
  assign w870[3] = |(datain[299:296] ^ 9);
  assign w870[4] = |(datain[295:292] ^ 12);
  assign w870[5] = |(datain[291:288] ^ 0);
  assign w870[6] = |(datain[287:284] ^ 12);
  assign w870[7] = |(datain[283:280] ^ 13);
  assign w870[8] = |(datain[279:276] ^ 2);
  assign w870[9] = |(datain[275:272] ^ 15);
  assign w870[10] = |(datain[271:268] ^ 14);
  assign w870[11] = |(datain[267:264] ^ 11);
  assign w870[12] = |(datain[263:260] ^ 0);
  assign w870[13] = |(datain[259:256] ^ 0);
  assign w870[14] = |(datain[255:252] ^ 0);
  assign w870[15] = |(datain[251:248] ^ 14);
  assign w870[16] = |(datain[247:244] ^ 1);
  assign w870[17] = |(datain[243:240] ^ 15);
  assign w870[18] = |(datain[239:236] ^ 12);
  assign w870[19] = |(datain[235:232] ^ 6);
  assign w870[20] = |(datain[231:228] ^ 0);
  assign w870[21] = |(datain[227:224] ^ 6);
  assign w870[22] = |(datain[223:220] ^ 14);
  assign w870[23] = |(datain[219:216] ^ 8);
  assign w870[24] = |(datain[215:212] ^ 0);
  assign w870[25] = |(datain[211:208] ^ 10);
  assign w870[26] = |(datain[207:204] ^ 0);
  assign w870[27] = |(datain[203:200] ^ 0);
  assign w870[28] = |(datain[199:196] ^ 14);
  assign w870[29] = |(datain[195:192] ^ 8);
  assign w870[30] = |(datain[191:188] ^ 13);
  assign w870[31] = |(datain[187:184] ^ 8);
  assign w870[32] = |(datain[183:180] ^ 0);
  assign w870[33] = |(datain[179:176] ^ 0);
  assign w870[34] = |(datain[175:172] ^ 11);
  assign w870[35] = |(datain[171:168] ^ 8);
  assign w870[36] = |(datain[167:164] ^ 0);
  assign w870[37] = |(datain[163:160] ^ 0);
  assign w870[38] = |(datain[159:156] ^ 1);
  assign w870[39] = |(datain[155:152] ^ 2);
  assign w870[40] = |(datain[151:148] ^ 12);
  assign w870[41] = |(datain[147:144] ^ 13);
  assign w870[42] = |(datain[143:140] ^ 2);
  assign w870[43] = |(datain[139:136] ^ 15);
  assign w870[44] = |(datain[135:132] ^ 15);
  assign w870[45] = |(datain[131:128] ^ 14);
  assign w870[46] = |(datain[127:124] ^ 12);
  assign w870[47] = |(datain[123:120] ^ 0);
  assign w870[48] = |(datain[119:116] ^ 7);
  assign w870[49] = |(datain[115:112] ^ 5);
  assign w870[50] = |(datain[111:108] ^ 0);
  assign w870[51] = |(datain[107:104] ^ 8);
  assign w870[52] = |(datain[103:100] ^ 11);
  assign w870[53] = |(datain[99:96] ^ 4);
  assign w870[54] = |(datain[95:92] ^ 3);
  assign w870[55] = |(datain[91:88] ^ 0);
  assign w870[56] = |(datain[87:84] ^ 12);
  assign w870[57] = |(datain[83:80] ^ 13);
  assign w870[58] = |(datain[79:76] ^ 2);
  assign w870[59] = |(datain[75:72] ^ 1);
  assign w870[60] = |(datain[71:68] ^ 3);
  assign w870[61] = |(datain[67:64] ^ 12);
  assign w870[62] = |(datain[63:60] ^ 0);
  assign w870[63] = |(datain[59:56] ^ 3);
  assign comp[870] = ~(|w870);
  wire [74-1:0] w871;
  assign w871[0] = |(datain[311:308] ^ 11);
  assign w871[1] = |(datain[307:304] ^ 10);
  assign w871[2] = |(datain[303:300] ^ 15);
  assign w871[3] = |(datain[299:296] ^ 10);
  assign w871[4] = |(datain[295:292] ^ 0);
  assign w871[5] = |(datain[291:288] ^ 10);
  assign w871[6] = |(datain[287:284] ^ 11);
  assign w871[7] = |(datain[283:280] ^ 8);
  assign w871[8] = |(datain[279:276] ^ 4);
  assign w871[9] = |(datain[275:272] ^ 0);
  assign w871[10] = |(datain[271:268] ^ 0);
  assign w871[11] = |(datain[267:264] ^ 0);
  assign w871[12] = |(datain[263:260] ^ 8);
  assign w871[13] = |(datain[259:256] ^ 6);
  assign w871[14] = |(datain[255:252] ^ 14);
  assign w871[15] = |(datain[251:248] ^ 0);
  assign w871[16] = |(datain[247:244] ^ 14);
  assign w871[17] = |(datain[243:240] ^ 8);
  assign w871[18] = |(datain[239:236] ^ 10);
  assign w871[19] = |(datain[235:232] ^ 13);
  assign w871[20] = |(datain[231:228] ^ 0);
  assign w871[21] = |(datain[227:224] ^ 1);
  assign w871[22] = |(datain[223:220] ^ 11);
  assign w871[23] = |(datain[219:216] ^ 8);
  assign w871[24] = |(datain[215:212] ^ 4);
  assign w871[25] = |(datain[211:208] ^ 2);
  assign w871[26] = |(datain[207:204] ^ 0);
  assign w871[27] = |(datain[203:200] ^ 0);
  assign w871[28] = |(datain[199:196] ^ 8);
  assign w871[29] = |(datain[195:192] ^ 6);
  assign w871[30] = |(datain[191:188] ^ 14);
  assign w871[31] = |(datain[187:184] ^ 0);
  assign w871[32] = |(datain[183:180] ^ 11);
  assign w871[33] = |(datain[179:176] ^ 10);
  assign w871[34] = |(datain[175:172] ^ 2);
  assign w871[35] = |(datain[171:168] ^ 6);
  assign w871[36] = |(datain[167:164] ^ 0);
  assign w871[37] = |(datain[163:160] ^ 0);
  assign w871[38] = |(datain[159:156] ^ 3);
  assign w871[39] = |(datain[155:152] ^ 3);
  assign w871[40] = |(datain[151:148] ^ 12);
  assign w871[41] = |(datain[147:144] ^ 9);
  assign w871[42] = |(datain[143:140] ^ 14);
  assign w871[43] = |(datain[139:136] ^ 8);
  assign w871[44] = |(datain[135:132] ^ 10);
  assign w871[45] = |(datain[131:128] ^ 0);
  assign w871[46] = |(datain[127:124] ^ 0);
  assign w871[47] = |(datain[123:120] ^ 1);
  assign w871[48] = |(datain[119:116] ^ 11);
  assign w871[49] = |(datain[115:112] ^ 8);
  assign w871[50] = |(datain[111:108] ^ 4);
  assign w871[51] = |(datain[107:104] ^ 2);
  assign w871[52] = |(datain[103:100] ^ 0);
  assign w871[53] = |(datain[99:96] ^ 0);
  assign w871[54] = |(datain[95:92] ^ 8);
  assign w871[55] = |(datain[91:88] ^ 6);
  assign w871[56] = |(datain[87:84] ^ 14);
  assign w871[57] = |(datain[83:80] ^ 0);
  assign w871[58] = |(datain[79:76] ^ 11);
  assign w871[59] = |(datain[75:72] ^ 10);
  assign w871[60] = |(datain[71:68] ^ 0);
  assign w871[61] = |(datain[67:64] ^ 6);
  assign w871[62] = |(datain[63:60] ^ 0);
  assign w871[63] = |(datain[59:56] ^ 2);
  assign w871[64] = |(datain[55:52] ^ 3);
  assign w871[65] = |(datain[51:48] ^ 3);
  assign w871[66] = |(datain[47:44] ^ 12);
  assign w871[67] = |(datain[43:40] ^ 9);
  assign w871[68] = |(datain[39:36] ^ 14);
  assign w871[69] = |(datain[35:32] ^ 8);
  assign w871[70] = |(datain[31:28] ^ 9);
  assign w871[71] = |(datain[27:24] ^ 3);
  assign w871[72] = |(datain[23:20] ^ 0);
  assign w871[73] = |(datain[19:16] ^ 1);
  assign comp[871] = ~(|w871);
  wire [72-1:0] w872;
  assign w872[0] = |(datain[311:308] ^ 0);
  assign w872[1] = |(datain[307:304] ^ 2);
  assign w872[2] = |(datain[303:300] ^ 9);
  assign w872[3] = |(datain[299:296] ^ 0);
  assign w872[4] = |(datain[295:292] ^ 11);
  assign w872[5] = |(datain[291:288] ^ 4);
  assign w872[6] = |(datain[287:284] ^ 4);
  assign w872[7] = |(datain[283:280] ^ 0);
  assign w872[8] = |(datain[279:276] ^ 12);
  assign w872[9] = |(datain[275:272] ^ 13);
  assign w872[10] = |(datain[271:268] ^ 2);
  assign w872[11] = |(datain[267:264] ^ 1);
  assign w872[12] = |(datain[263:260] ^ 11);
  assign w872[13] = |(datain[259:256] ^ 8);
  assign w872[14] = |(datain[255:252] ^ 0);
  assign w872[15] = |(datain[251:248] ^ 0);
  assign w872[16] = |(datain[247:244] ^ 4);
  assign w872[17] = |(datain[243:240] ^ 2);
  assign w872[18] = |(datain[239:236] ^ 3);
  assign w872[19] = |(datain[235:232] ^ 3);
  assign w872[20] = |(datain[231:228] ^ 12);
  assign w872[21] = |(datain[227:224] ^ 9);
  assign w872[22] = |(datain[223:220] ^ 3);
  assign w872[23] = |(datain[219:216] ^ 3);
  assign w872[24] = |(datain[215:212] ^ 13);
  assign w872[25] = |(datain[211:208] ^ 2);
  assign w872[26] = |(datain[207:204] ^ 12);
  assign w872[27] = |(datain[203:200] ^ 13);
  assign w872[28] = |(datain[199:196] ^ 2);
  assign w872[29] = |(datain[195:192] ^ 1);
  assign w872[30] = |(datain[191:188] ^ 8);
  assign w872[31] = |(datain[187:184] ^ 1);
  assign w872[32] = |(datain[183:180] ^ 12);
  assign w872[33] = |(datain[179:176] ^ 7);
  assign w872[34] = |(datain[175:172] ^ 7);
  assign w872[35] = |(datain[171:168] ^ 3);
  assign w872[36] = |(datain[167:164] ^ 0);
  assign w872[37] = |(datain[163:160] ^ 2);
  assign w872[38] = |(datain[159:156] ^ 12);
  assign w872[39] = |(datain[155:152] ^ 6);
  assign w872[40] = |(datain[151:148] ^ 0);
  assign w872[41] = |(datain[147:144] ^ 5);
  assign w872[42] = |(datain[143:140] ^ 0);
  assign w872[43] = |(datain[139:136] ^ 3);
  assign w872[44] = |(datain[135:132] ^ 12);
  assign w872[45] = |(datain[131:128] ^ 6);
  assign w872[46] = |(datain[127:124] ^ 4);
  assign w872[47] = |(datain[123:120] ^ 5);
  assign w872[48] = |(datain[119:116] ^ 0);
  assign w872[49] = |(datain[115:112] ^ 1);
  assign w872[50] = |(datain[111:108] ^ 0);
  assign w872[51] = |(datain[107:104] ^ 1);
  assign w872[52] = |(datain[103:100] ^ 8);
  assign w872[53] = |(datain[99:96] ^ 11);
  assign w872[54] = |(datain[95:92] ^ 4);
  assign w872[55] = |(datain[91:88] ^ 5);
  assign w872[56] = |(datain[87:84] ^ 1);
  assign w872[57] = |(datain[83:80] ^ 15);
  assign w872[58] = |(datain[79:76] ^ 12);
  assign w872[59] = |(datain[75:72] ^ 6);
  assign w872[60] = |(datain[71:68] ^ 4);
  assign w872[61] = |(datain[67:64] ^ 5);
  assign w872[62] = |(datain[63:60] ^ 0);
  assign w872[63] = |(datain[59:56] ^ 2);
  assign w872[64] = |(datain[55:52] ^ 14);
  assign w872[65] = |(datain[51:48] ^ 9);
  assign w872[66] = |(datain[47:44] ^ 2);
  assign w872[67] = |(datain[43:40] ^ 13);
  assign w872[68] = |(datain[39:36] ^ 0);
  assign w872[69] = |(datain[35:32] ^ 5);
  assign w872[70] = |(datain[31:28] ^ 0);
  assign w872[71] = |(datain[27:24] ^ 0);
  assign comp[872] = ~(|w872);
  wire [76-1:0] w873;
  assign w873[0] = |(datain[311:308] ^ 15);
  assign w873[1] = |(datain[307:304] ^ 0);
  assign w873[2] = |(datain[303:300] ^ 3);
  assign w873[3] = |(datain[299:296] ^ 13);
  assign w873[4] = |(datain[295:292] ^ 0);
  assign w873[5] = |(datain[291:288] ^ 0);
  assign w873[6] = |(datain[287:284] ^ 15);
  assign w873[7] = |(datain[283:280] ^ 0);
  assign w873[8] = |(datain[279:276] ^ 7);
  assign w873[9] = |(datain[275:272] ^ 5);
  assign w873[10] = |(datain[271:268] ^ 0);
  assign w873[11] = |(datain[267:264] ^ 3);
  assign w873[12] = |(datain[263:260] ^ 14);
  assign w873[13] = |(datain[259:256] ^ 9);
  assign w873[14] = |(datain[255:252] ^ 3);
  assign w873[15] = |(datain[251:248] ^ 3);
  assign w873[16] = |(datain[247:244] ^ 0);
  assign w873[17] = |(datain[243:240] ^ 0);
  assign w873[18] = |(datain[239:236] ^ 8);
  assign w873[19] = |(datain[235:232] ^ 11);
  assign w873[20] = |(datain[231:228] ^ 13);
  assign w873[21] = |(datain[227:224] ^ 5);
  assign w873[22] = |(datain[223:220] ^ 11);
  assign w873[23] = |(datain[219:216] ^ 9);
  assign w873[24] = |(datain[215:212] ^ 7);
  assign w873[25] = |(datain[211:208] ^ 1);
  assign w873[26] = |(datain[207:204] ^ 0);
  assign w873[27] = |(datain[203:200] ^ 2);
  assign w873[28] = |(datain[199:196] ^ 11);
  assign w873[29] = |(datain[195:192] ^ 4);
  assign w873[30] = |(datain[191:188] ^ 4);
  assign w873[31] = |(datain[187:184] ^ 0);
  assign w873[32] = |(datain[183:180] ^ 12);
  assign w873[33] = |(datain[179:176] ^ 13);
  assign w873[34] = |(datain[175:172] ^ 2);
  assign w873[35] = |(datain[171:168] ^ 1);
  assign w873[36] = |(datain[167:164] ^ 11);
  assign w873[37] = |(datain[163:160] ^ 8);
  assign w873[38] = |(datain[159:156] ^ 0);
  assign w873[39] = |(datain[155:152] ^ 0);
  assign w873[40] = |(datain[151:148] ^ 4);
  assign w873[41] = |(datain[147:144] ^ 2);
  assign w873[42] = |(datain[143:140] ^ 3);
  assign w873[43] = |(datain[139:136] ^ 3);
  assign w873[44] = |(datain[135:132] ^ 12);
  assign w873[45] = |(datain[131:128] ^ 9);
  assign w873[46] = |(datain[127:124] ^ 3);
  assign w873[47] = |(datain[123:120] ^ 3);
  assign w873[48] = |(datain[119:116] ^ 13);
  assign w873[49] = |(datain[115:112] ^ 2);
  assign w873[50] = |(datain[111:108] ^ 12);
  assign w873[51] = |(datain[107:104] ^ 13);
  assign w873[52] = |(datain[103:100] ^ 2);
  assign w873[53] = |(datain[99:96] ^ 1);
  assign w873[54] = |(datain[95:92] ^ 8);
  assign w873[55] = |(datain[91:88] ^ 1);
  assign w873[56] = |(datain[87:84] ^ 12);
  assign w873[57] = |(datain[83:80] ^ 7);
  assign w873[58] = |(datain[79:76] ^ 7);
  assign w873[59] = |(datain[75:72] ^ 1);
  assign w873[60] = |(datain[71:68] ^ 0);
  assign w873[61] = |(datain[67:64] ^ 2);
  assign w873[62] = |(datain[63:60] ^ 12);
  assign w873[63] = |(datain[59:56] ^ 6);
  assign w873[64] = |(datain[55:52] ^ 0);
  assign w873[65] = |(datain[51:48] ^ 5);
  assign w873[66] = |(datain[47:44] ^ 0);
  assign w873[67] = |(datain[43:40] ^ 3);
  assign w873[68] = |(datain[39:36] ^ 12);
  assign w873[69] = |(datain[35:32] ^ 6);
  assign w873[70] = |(datain[31:28] ^ 4);
  assign w873[71] = |(datain[27:24] ^ 5);
  assign w873[72] = |(datain[23:20] ^ 0);
  assign w873[73] = |(datain[19:16] ^ 1);
  assign w873[74] = |(datain[15:12] ^ 0);
  assign w873[75] = |(datain[11:8] ^ 1);
  assign comp[873] = ~(|w873);
  wire [42-1:0] w874;
  assign w874[0] = |(datain[311:308] ^ 0);
  assign w874[1] = |(datain[307:304] ^ 3);
  assign w874[2] = |(datain[303:300] ^ 13);
  assign w874[3] = |(datain[299:296] ^ 6);
  assign w874[4] = |(datain[295:292] ^ 12);
  assign w874[5] = |(datain[291:288] ^ 13);
  assign w874[6] = |(datain[287:284] ^ 2);
  assign w874[7] = |(datain[283:280] ^ 1);
  assign w874[8] = |(datain[279:276] ^ 1);
  assign w874[9] = |(datain[275:272] ^ 14);
  assign w874[10] = |(datain[271:268] ^ 0);
  assign w874[11] = |(datain[267:264] ^ 7);
  assign w874[12] = |(datain[263:260] ^ 0);
  assign w874[13] = |(datain[259:256] ^ 6);
  assign w874[14] = |(datain[255:252] ^ 11);
  assign w874[15] = |(datain[251:248] ^ 4);
  assign w874[16] = |(datain[247:244] ^ 2);
  assign w874[17] = |(datain[243:240] ^ 15);
  assign w874[18] = |(datain[239:236] ^ 12);
  assign w874[19] = |(datain[235:232] ^ 13);
  assign w874[20] = |(datain[231:228] ^ 2);
  assign w874[21] = |(datain[227:224] ^ 1);
  assign w874[22] = |(datain[223:220] ^ 8);
  assign w874[23] = |(datain[219:216] ^ 12);
  assign w874[24] = |(datain[215:212] ^ 4);
  assign w874[25] = |(datain[211:208] ^ 4);
  assign w874[26] = |(datain[207:204] ^ 4);
  assign w874[27] = |(datain[203:200] ^ 10);
  assign w874[28] = |(datain[199:196] ^ 8);
  assign w874[29] = |(datain[195:192] ^ 9);
  assign w874[30] = |(datain[191:188] ^ 5);
  assign w874[31] = |(datain[187:184] ^ 12);
  assign w874[32] = |(datain[183:180] ^ 4);
  assign w874[33] = |(datain[179:176] ^ 12);
  assign w874[34] = |(datain[175:172] ^ 0);
  assign w874[35] = |(datain[171:168] ^ 7);
  assign w874[36] = |(datain[167:164] ^ 11);
  assign w874[37] = |(datain[163:160] ^ 4);
  assign w874[38] = |(datain[159:156] ^ 1);
  assign w874[39] = |(datain[155:152] ^ 10);
  assign w874[40] = |(datain[151:148] ^ 11);
  assign w874[41] = |(datain[147:144] ^ 10);
  assign comp[874] = ~(|w874);
  wire [30-1:0] w875;
  assign w875[0] = |(datain[311:308] ^ 11);
  assign w875[1] = |(datain[307:304] ^ 10);
  assign w875[2] = |(datain[303:300] ^ 12);
  assign w875[3] = |(datain[299:296] ^ 12);
  assign w875[4] = |(datain[295:292] ^ 0);
  assign w875[5] = |(datain[291:288] ^ 2);
  assign w875[6] = |(datain[287:284] ^ 11);
  assign w875[7] = |(datain[283:280] ^ 4);
  assign w875[8] = |(datain[279:276] ^ 0);
  assign w875[9] = |(datain[275:272] ^ 9);
  assign w875[10] = |(datain[271:268] ^ 12);
  assign w875[11] = |(datain[267:264] ^ 13);
  assign w875[12] = |(datain[263:260] ^ 2);
  assign w875[13] = |(datain[259:256] ^ 1);
  assign w875[14] = |(datain[255:252] ^ 11);
  assign w875[15] = |(datain[251:248] ^ 4);
  assign w875[16] = |(datain[247:244] ^ 4);
  assign w875[17] = |(datain[243:240] ^ 12);
  assign w875[18] = |(datain[239:236] ^ 12);
  assign w875[19] = |(datain[235:232] ^ 13);
  assign w875[20] = |(datain[231:228] ^ 2);
  assign w875[21] = |(datain[227:224] ^ 1);
  assign w875[22] = |(datain[223:220] ^ 11);
  assign w875[23] = |(datain[219:216] ^ 10);
  assign w875[24] = |(datain[215:212] ^ 0);
  assign w875[25] = |(datain[211:208] ^ 0);
  assign w875[26] = |(datain[207:204] ^ 0);
  assign w875[27] = |(datain[203:200] ^ 3);
  assign w875[28] = |(datain[199:196] ^ 11);
  assign w875[29] = |(datain[195:192] ^ 4);
  assign comp[875] = ~(|w875);
  wire [44-1:0] w876;
  assign w876[0] = |(datain[311:308] ^ 3);
  assign w876[1] = |(datain[307:304] ^ 14);
  assign w876[2] = |(datain[303:300] ^ 0);
  assign w876[3] = |(datain[299:296] ^ 0);
  assign w876[4] = |(datain[295:292] ^ 11);
  assign w876[5] = |(datain[291:288] ^ 9);
  assign w876[6] = |(datain[287:284] ^ 14);
  assign w876[7] = |(datain[283:280] ^ 13);
  assign w876[8] = |(datain[279:276] ^ 0);
  assign w876[9] = |(datain[275:272] ^ 2);
  assign w876[10] = |(datain[271:268] ^ 8);
  assign w876[11] = |(datain[267:264] ^ 10);
  assign w876[12] = |(datain[263:260] ^ 0);
  assign w876[13] = |(datain[259:256] ^ 7);
  assign w876[14] = |(datain[255:252] ^ 14);
  assign w876[15] = |(datain[251:248] ^ 8);
  assign w876[16] = |(datain[247:244] ^ 0);
  assign w876[17] = |(datain[243:240] ^ 8);
  assign w876[18] = |(datain[239:236] ^ 0);
  assign w876[19] = |(datain[235:232] ^ 0);
  assign w876[20] = |(datain[231:228] ^ 8);
  assign w876[21] = |(datain[227:224] ^ 8);
  assign w876[22] = |(datain[223:220] ^ 0);
  assign w876[23] = |(datain[219:216] ^ 7);
  assign w876[24] = |(datain[215:212] ^ 4);
  assign w876[25] = |(datain[211:208] ^ 3);
  assign w876[26] = |(datain[207:204] ^ 14);
  assign w876[27] = |(datain[203:200] ^ 2);
  assign w876[28] = |(datain[199:196] ^ 15);
  assign w876[29] = |(datain[195:192] ^ 6);
  assign w876[30] = |(datain[191:188] ^ 1);
  assign w876[31] = |(datain[187:184] ^ 15);
  assign w876[32] = |(datain[183:180] ^ 14);
  assign w876[33] = |(datain[179:176] ^ 11);
  assign w876[34] = |(datain[175:172] ^ 1);
  assign w876[35] = |(datain[171:168] ^ 2);
  assign w876[36] = |(datain[167:164] ^ 5);
  assign w876[37] = |(datain[163:160] ^ 0);
  assign w876[38] = |(datain[159:156] ^ 5);
  assign w876[39] = |(datain[155:152] ^ 3);
  assign w876[40] = |(datain[151:148] ^ 5);
  assign w876[41] = |(datain[147:144] ^ 1);
  assign w876[42] = |(datain[143:140] ^ 11);
  assign w876[43] = |(datain[139:136] ^ 8);
  assign comp[876] = ~(|w876);
  wire [46-1:0] w877;
  assign w877[0] = |(datain[311:308] ^ 12);
  assign w877[1] = |(datain[307:304] ^ 3);
  assign w877[2] = |(datain[303:300] ^ 3);
  assign w877[3] = |(datain[299:296] ^ 14);
  assign w877[4] = |(datain[295:292] ^ 0);
  assign w877[5] = |(datain[291:288] ^ 0);
  assign w877[6] = |(datain[287:284] ^ 11);
  assign w877[7] = |(datain[283:280] ^ 9);
  assign w877[8] = |(datain[279:276] ^ 14);
  assign w877[9] = |(datain[275:272] ^ 12);
  assign w877[10] = |(datain[271:268] ^ 0);
  assign w877[11] = |(datain[267:264] ^ 2);
  assign w877[12] = |(datain[263:260] ^ 8);
  assign w877[13] = |(datain[259:256] ^ 10);
  assign w877[14] = |(datain[255:252] ^ 0);
  assign w877[15] = |(datain[251:248] ^ 7);
  assign w877[16] = |(datain[247:244] ^ 14);
  assign w877[17] = |(datain[243:240] ^ 8);
  assign w877[18] = |(datain[239:236] ^ 0);
  assign w877[19] = |(datain[235:232] ^ 8);
  assign w877[20] = |(datain[231:228] ^ 0);
  assign w877[21] = |(datain[227:224] ^ 0);
  assign w877[22] = |(datain[223:220] ^ 8);
  assign w877[23] = |(datain[219:216] ^ 8);
  assign w877[24] = |(datain[215:212] ^ 0);
  assign w877[25] = |(datain[211:208] ^ 7);
  assign w877[26] = |(datain[207:204] ^ 4);
  assign w877[27] = |(datain[203:200] ^ 3);
  assign w877[28] = |(datain[199:196] ^ 14);
  assign w877[29] = |(datain[195:192] ^ 2);
  assign w877[30] = |(datain[191:188] ^ 15);
  assign w877[31] = |(datain[187:184] ^ 6);
  assign w877[32] = |(datain[183:180] ^ 1);
  assign w877[33] = |(datain[179:176] ^ 15);
  assign w877[34] = |(datain[175:172] ^ 14);
  assign w877[35] = |(datain[171:168] ^ 11);
  assign w877[36] = |(datain[167:164] ^ 1);
  assign w877[37] = |(datain[163:160] ^ 2);
  assign w877[38] = |(datain[159:156] ^ 5);
  assign w877[39] = |(datain[155:152] ^ 0);
  assign w877[40] = |(datain[151:148] ^ 5);
  assign w877[41] = |(datain[147:144] ^ 3);
  assign w877[42] = |(datain[143:140] ^ 5);
  assign w877[43] = |(datain[139:136] ^ 1);
  assign w877[44] = |(datain[135:132] ^ 11);
  assign w877[45] = |(datain[131:128] ^ 8);
  assign comp[877] = ~(|w877);
  wire [44-1:0] w878;
  assign w878[0] = |(datain[311:308] ^ 8);
  assign w878[1] = |(datain[307:304] ^ 14);
  assign w878[2] = |(datain[303:300] ^ 13);
  assign w878[3] = |(datain[299:296] ^ 9);
  assign w878[4] = |(datain[295:292] ^ 11);
  assign w878[5] = |(datain[291:288] ^ 14);
  assign w878[6] = |(datain[287:284] ^ 8);
  assign w878[7] = |(datain[283:280] ^ 4);
  assign w878[8] = |(datain[279:276] ^ 0);
  assign w878[9] = |(datain[275:272] ^ 0);
  assign w878[10] = |(datain[271:268] ^ 11);
  assign w878[11] = |(datain[267:264] ^ 15);
  assign w878[12] = |(datain[263:260] ^ 0);
  assign w878[13] = |(datain[259:256] ^ 8);
  assign w878[14] = |(datain[255:252] ^ 0);
  assign w878[15] = |(datain[251:248] ^ 3);
  assign w878[16] = |(datain[247:244] ^ 11);
  assign w878[17] = |(datain[243:240] ^ 10);
  assign w878[18] = |(datain[239:236] ^ 5);
  assign w878[19] = |(datain[235:232] ^ 11);
  assign w878[20] = |(datain[231:228] ^ 0);
  assign w878[21] = |(datain[227:224] ^ 1);
  assign w878[22] = |(datain[223:220] ^ 10);
  assign w878[23] = |(datain[219:216] ^ 13);
  assign w878[24] = |(datain[215:212] ^ 3);
  assign w878[25] = |(datain[211:208] ^ 11);
  assign w878[26] = |(datain[207:204] ^ 12);
  assign w878[27] = |(datain[203:200] ^ 2);
  assign w878[28] = |(datain[199:196] ^ 7);
  assign w878[29] = |(datain[195:192] ^ 4);
  assign w878[30] = |(datain[191:188] ^ 0);
  assign w878[31] = |(datain[187:184] ^ 11);
  assign w878[32] = |(datain[183:180] ^ 10);
  assign w878[33] = |(datain[179:176] ^ 11);
  assign w878[34] = |(datain[175:172] ^ 10);
  assign w878[35] = |(datain[171:168] ^ 5);
  assign w878[36] = |(datain[167:164] ^ 0);
  assign w878[37] = |(datain[163:160] ^ 6);
  assign w878[38] = |(datain[159:156] ^ 1);
  assign w878[39] = |(datain[155:152] ^ 15);
  assign w878[40] = |(datain[151:148] ^ 11);
  assign w878[41] = |(datain[147:144] ^ 8);
  assign w878[42] = |(datain[143:140] ^ 2);
  assign w878[43] = |(datain[139:136] ^ 1);
  assign comp[878] = ~(|w878);
  wire [50-1:0] w879;
  assign w879[0] = |(datain[311:308] ^ 11);
  assign w879[1] = |(datain[307:304] ^ 4);
  assign w879[2] = |(datain[303:300] ^ 0);
  assign w879[3] = |(datain[299:296] ^ 8);
  assign w879[4] = |(datain[295:292] ^ 11);
  assign w879[5] = |(datain[291:288] ^ 2);
  assign w879[6] = |(datain[287:284] ^ 14);
  assign w879[7] = |(datain[283:280] ^ 0);
  assign w879[8] = |(datain[279:276] ^ 12);
  assign w879[9] = |(datain[275:272] ^ 13);
  assign w879[10] = |(datain[271:268] ^ 1);
  assign w879[11] = |(datain[267:264] ^ 3);
  assign w879[12] = |(datain[263:260] ^ 8);
  assign w879[13] = |(datain[259:256] ^ 0);
  assign w879[14] = |(datain[255:252] ^ 12);
  assign w879[15] = |(datain[251:248] ^ 4);
  assign w879[16] = |(datain[247:244] ^ 0);
  assign w879[17] = |(datain[243:240] ^ 11);
  assign w879[18] = |(datain[239:236] ^ 11);
  assign w879[19] = |(datain[235:232] ^ 9);
  assign w879[20] = |(datain[231:228] ^ 7);
  assign w879[21] = |(datain[227:224] ^ 14);
  assign w879[22] = |(datain[223:220] ^ 0);
  assign w879[23] = |(datain[219:216] ^ 1);
  assign w879[24] = |(datain[215:212] ^ 2);
  assign w879[25] = |(datain[211:208] ^ 14);
  assign w879[26] = |(datain[207:204] ^ 8);
  assign w879[27] = |(datain[203:200] ^ 10);
  assign w879[28] = |(datain[199:196] ^ 0);
  assign w879[29] = |(datain[195:192] ^ 4);
  assign w879[30] = |(datain[191:188] ^ 3);
  assign w879[31] = |(datain[187:184] ^ 2);
  assign w879[32] = |(datain[183:180] ^ 12);
  assign w879[33] = |(datain[179:176] ^ 4);
  assign w879[34] = |(datain[175:172] ^ 2);
  assign w879[35] = |(datain[171:168] ^ 14);
  assign w879[36] = |(datain[167:164] ^ 8);
  assign w879[37] = |(datain[163:160] ^ 8);
  assign w879[38] = |(datain[159:156] ^ 0);
  assign w879[39] = |(datain[155:152] ^ 4);
  assign w879[40] = |(datain[151:148] ^ 4);
  assign w879[41] = |(datain[147:144] ^ 6);
  assign w879[42] = |(datain[143:140] ^ 14);
  assign w879[43] = |(datain[139:136] ^ 2);
  assign w879[44] = |(datain[135:132] ^ 15);
  assign w879[45] = |(datain[131:128] ^ 5);
  assign w879[46] = |(datain[127:124] ^ 6);
  assign w879[47] = |(datain[123:120] ^ 1);
  assign w879[48] = |(datain[119:116] ^ 12);
  assign w879[49] = |(datain[115:112] ^ 3);
  assign comp[879] = ~(|w879);
  wire [40-1:0] w880;
  assign w880[0] = |(datain[311:308] ^ 14);
  assign w880[1] = |(datain[307:304] ^ 2);
  assign w880[2] = |(datain[303:300] ^ 15);
  assign w880[3] = |(datain[299:296] ^ 10);
  assign w880[4] = |(datain[295:292] ^ 5);
  assign w880[5] = |(datain[291:288] ^ 11);
  assign w880[6] = |(datain[287:284] ^ 5);
  assign w880[7] = |(datain[283:280] ^ 9);
  assign w880[8] = |(datain[279:276] ^ 5);
  assign w880[9] = |(datain[275:272] ^ 8);
  assign w880[10] = |(datain[271:268] ^ 5);
  assign w880[11] = |(datain[267:264] ^ 14);
  assign w880[12] = |(datain[263:260] ^ 12);
  assign w880[13] = |(datain[259:256] ^ 3);
  assign w880[14] = |(datain[255:252] ^ 14);
  assign w880[15] = |(datain[251:248] ^ 8);
  assign w880[16] = |(datain[247:244] ^ 13);
  assign w880[17] = |(datain[243:240] ^ 12);
  assign w880[18] = |(datain[239:236] ^ 15);
  assign w880[19] = |(datain[235:232] ^ 15);
  assign w880[20] = |(datain[231:228] ^ 8);
  assign w880[21] = |(datain[227:224] ^ 9);
  assign w880[22] = |(datain[223:220] ^ 8);
  assign w880[23] = |(datain[219:216] ^ 4);
  assign w880[24] = |(datain[215:212] ^ 14);
  assign w880[25] = |(datain[211:208] ^ 4);
  assign w880[26] = |(datain[207:204] ^ 0);
  assign w880[27] = |(datain[203:200] ^ 2);
  assign w880[28] = |(datain[199:196] ^ 8);
  assign w880[29] = |(datain[195:192] ^ 13);
  assign w880[30] = |(datain[191:188] ^ 9);
  assign w880[31] = |(datain[187:184] ^ 4);
  assign w880[32] = |(datain[183:180] ^ 0);
  assign w880[33] = |(datain[179:176] ^ 5);
  assign w880[34] = |(datain[175:172] ^ 0);
  assign w880[35] = |(datain[171:168] ^ 1);
  assign w880[36] = |(datain[167:164] ^ 11);
  assign w880[37] = |(datain[163:160] ^ 4);
  assign w880[38] = |(datain[159:156] ^ 4);
  assign w880[39] = |(datain[155:152] ^ 0);
  assign comp[880] = ~(|w880);
  wire [32-1:0] w881;
  assign w881[0] = |(datain[311:308] ^ 11);
  assign w881[1] = |(datain[307:304] ^ 8);
  assign w881[2] = |(datain[303:300] ^ 0);
  assign w881[3] = |(datain[299:296] ^ 0);
  assign w881[4] = |(datain[295:292] ^ 1);
  assign w881[5] = |(datain[291:288] ^ 10);
  assign w881[6] = |(datain[287:284] ^ 12);
  assign w881[7] = |(datain[283:280] ^ 13);
  assign w881[8] = |(datain[279:276] ^ 2);
  assign w881[9] = |(datain[275:272] ^ 1);
  assign w881[10] = |(datain[271:268] ^ 5);
  assign w881[11] = |(datain[267:264] ^ 14);
  assign w881[12] = |(datain[263:260] ^ 8);
  assign w881[13] = |(datain[259:256] ^ 11);
  assign w881[14] = |(datain[255:252] ^ 1);
  assign w881[15] = |(datain[251:248] ^ 12);
  assign w881[16] = |(datain[247:244] ^ 11);
  assign w881[17] = |(datain[243:240] ^ 9);
  assign w881[18] = |(datain[239:236] ^ 0);
  assign w881[19] = |(datain[235:232] ^ 3);
  assign w881[20] = |(datain[231:228] ^ 0);
  assign w881[21] = |(datain[227:224] ^ 8);
  assign w881[22] = |(datain[223:220] ^ 11);
  assign w881[23] = |(datain[219:216] ^ 8);
  assign w881[24] = |(datain[215:212] ^ 0);
  assign w881[25] = |(datain[211:208] ^ 0);
  assign w881[26] = |(datain[207:204] ^ 4);
  assign w881[27] = |(datain[203:200] ^ 0);
  assign w881[28] = |(datain[199:196] ^ 12);
  assign w881[29] = |(datain[195:192] ^ 13);
  assign w881[30] = |(datain[191:188] ^ 2);
  assign w881[31] = |(datain[187:184] ^ 1);
  assign comp[881] = ~(|w881);
  wire [46-1:0] w882;
  assign w882[0] = |(datain[311:308] ^ 9);
  assign w882[1] = |(datain[307:304] ^ 13);
  assign w882[2] = |(datain[303:300] ^ 8);
  assign w882[3] = |(datain[299:296] ^ 1);
  assign w882[4] = |(datain[295:292] ^ 15);
  assign w882[5] = |(datain[291:288] ^ 9);
  assign w882[6] = |(datain[287:284] ^ 15);
  assign w882[7] = |(datain[283:280] ^ 14);
  assign w882[8] = |(datain[279:276] ^ 15);
  assign w882[9] = |(datain[275:272] ^ 10);
  assign w882[10] = |(datain[271:268] ^ 7);
  assign w882[11] = |(datain[267:264] ^ 5);
  assign w882[12] = |(datain[263:260] ^ 1);
  assign w882[13] = |(datain[259:256] ^ 0);
  assign w882[14] = |(datain[255:252] ^ 8);
  assign w882[15] = |(datain[251:248] ^ 1);
  assign w882[16] = |(datain[247:244] ^ 15);
  assign w882[17] = |(datain[243:240] ^ 10);
  assign w882[18] = |(datain[239:236] ^ 15);
  assign w882[19] = |(datain[235:232] ^ 10);
  assign w882[20] = |(datain[231:228] ^ 15);
  assign w882[21] = |(datain[227:224] ^ 14);
  assign w882[22] = |(datain[223:220] ^ 7);
  assign w882[23] = |(datain[219:216] ^ 5);
  assign w882[24] = |(datain[215:212] ^ 0);
  assign w882[25] = |(datain[211:208] ^ 10);
  assign w882[26] = |(datain[207:204] ^ 15);
  assign w882[27] = |(datain[203:200] ^ 10);
  assign w882[28] = |(datain[199:196] ^ 9);
  assign w882[29] = |(datain[195:192] ^ 12);
  assign w882[30] = |(datain[191:188] ^ 2);
  assign w882[31] = |(datain[187:184] ^ 14);
  assign w882[32] = |(datain[183:180] ^ 15);
  assign w882[33] = |(datain[179:176] ^ 15);
  assign w882[34] = |(datain[175:172] ^ 1);
  assign w882[35] = |(datain[171:168] ^ 14);
  assign w882[36] = |(datain[167:164] ^ 9);
  assign w882[37] = |(datain[163:160] ^ 14);
  assign w882[38] = |(datain[159:156] ^ 0);
  assign w882[39] = |(datain[155:152] ^ 0);
  assign w882[40] = |(datain[151:148] ^ 11);
  assign w882[41] = |(datain[147:144] ^ 9);
  assign w882[42] = |(datain[143:140] ^ 14);
  assign w882[43] = |(datain[139:136] ^ 14);
  assign w882[44] = |(datain[135:132] ^ 14);
  assign w882[45] = |(datain[131:128] ^ 14);
  assign comp[882] = ~(|w882);
  wire [74-1:0] w883;
  assign w883[0] = |(datain[311:308] ^ 11);
  assign w883[1] = |(datain[307:304] ^ 15);
  assign w883[2] = |(datain[303:300] ^ 9);
  assign w883[3] = |(datain[299:296] ^ 14);
  assign w883[4] = |(datain[295:292] ^ 0);
  assign w883[5] = |(datain[291:288] ^ 0);
  assign w883[6] = |(datain[287:284] ^ 11);
  assign w883[7] = |(datain[283:280] ^ 0);
  assign w883[8] = |(datain[279:276] ^ 0);
  assign w883[9] = |(datain[275:272] ^ 0);
  assign w883[10] = |(datain[271:268] ^ 11);
  assign w883[11] = |(datain[267:264] ^ 9);
  assign w883[12] = |(datain[263:260] ^ 0);
  assign w883[13] = |(datain[259:256] ^ 12);
  assign w883[14] = |(datain[255:252] ^ 0);
  assign w883[15] = |(datain[251:248] ^ 0);
  assign w883[16] = |(datain[247:244] ^ 15);
  assign w883[17] = |(datain[243:240] ^ 2);
  assign w883[18] = |(datain[239:236] ^ 10);
  assign w883[19] = |(datain[235:232] ^ 14);
  assign w883[20] = |(datain[231:228] ^ 12);
  assign w883[21] = |(datain[227:224] ^ 6);
  assign w883[22] = |(datain[223:220] ^ 0);
  assign w883[23] = |(datain[219:216] ^ 5);
  assign w883[24] = |(datain[215:212] ^ 0);
  assign w883[25] = |(datain[211:208] ^ 0);
  assign w883[26] = |(datain[207:204] ^ 11);
  assign w883[27] = |(datain[203:200] ^ 4);
  assign w883[28] = |(datain[199:196] ^ 3);
  assign w883[29] = |(datain[195:192] ^ 13);
  assign w883[30] = |(datain[191:188] ^ 11);
  assign w883[31] = |(datain[187:184] ^ 0);
  assign w883[32] = |(datain[183:180] ^ 0);
  assign w883[33] = |(datain[179:176] ^ 1);
  assign w883[34] = |(datain[175:172] ^ 12);
  assign w883[35] = |(datain[171:168] ^ 13);
  assign w883[36] = |(datain[167:164] ^ 2);
  assign w883[37] = |(datain[163:160] ^ 1);
  assign w883[38] = |(datain[159:156] ^ 8);
  assign w883[39] = |(datain[155:152] ^ 9);
  assign w883[40] = |(datain[151:148] ^ 12);
  assign w883[41] = |(datain[147:144] ^ 3);
  assign w883[42] = |(datain[143:140] ^ 11);
  assign w883[43] = |(datain[139:136] ^ 4);
  assign w883[44] = |(datain[135:132] ^ 4);
  assign w883[45] = |(datain[131:128] ^ 0);
  assign w883[46] = |(datain[127:124] ^ 11);
  assign w883[47] = |(datain[123:120] ^ 10);
  assign w883[48] = |(datain[119:116] ^ 0);
  assign w883[49] = |(datain[115:112] ^ 0);
  assign w883[50] = |(datain[111:108] ^ 0);
  assign w883[51] = |(datain[107:104] ^ 1);
  assign w883[52] = |(datain[103:100] ^ 11);
  assign w883[53] = |(datain[99:96] ^ 9);
  assign w883[54] = |(datain[95:92] ^ 1);
  assign w883[55] = |(datain[91:88] ^ 12);
  assign w883[56] = |(datain[87:84] ^ 0);
  assign w883[57] = |(datain[83:80] ^ 1);
  assign w883[58] = |(datain[79:76] ^ 12);
  assign w883[59] = |(datain[75:72] ^ 13);
  assign w883[60] = |(datain[71:68] ^ 2);
  assign w883[61] = |(datain[67:64] ^ 1);
  assign w883[62] = |(datain[63:60] ^ 11);
  assign w883[63] = |(datain[59:56] ^ 4);
  assign w883[64] = |(datain[55:52] ^ 3);
  assign w883[65] = |(datain[51:48] ^ 14);
  assign w883[66] = |(datain[47:44] ^ 12);
  assign w883[67] = |(datain[43:40] ^ 13);
  assign w883[68] = |(datain[39:36] ^ 2);
  assign w883[69] = |(datain[35:32] ^ 1);
  assign w883[70] = |(datain[31:28] ^ 11);
  assign w883[71] = |(datain[27:24] ^ 4);
  assign w883[72] = |(datain[23:20] ^ 4);
  assign w883[73] = |(datain[19:16] ^ 14);
  assign comp[883] = ~(|w883);
  wire [46-1:0] w884;
  assign w884[0] = |(datain[311:308] ^ 12);
  assign w884[1] = |(datain[307:304] ^ 15);
  assign w884[2] = |(datain[303:300] ^ 14);
  assign w884[3] = |(datain[299:296] ^ 11);
  assign w884[4] = |(datain[295:292] ^ 0);
  assign w884[5] = |(datain[291:288] ^ 3);
  assign w884[6] = |(datain[287:284] ^ 9);
  assign w884[7] = |(datain[283:280] ^ 0);
  assign w884[8] = |(datain[279:276] ^ 15);
  assign w884[9] = |(datain[275:272] ^ 13);
  assign w884[10] = |(datain[271:268] ^ 13);
  assign w884[11] = |(datain[267:264] ^ 3);
  assign w884[12] = |(datain[263:260] ^ 8);
  assign w884[13] = |(datain[259:256] ^ 10);
  assign w884[14] = |(datain[255:252] ^ 10);
  assign w884[15] = |(datain[251:248] ^ 6);
  assign w884[16] = |(datain[247:244] ^ 4);
  assign w884[17] = |(datain[243:240] ^ 9);
  assign w884[18] = |(datain[239:236] ^ 0);
  assign w884[19] = |(datain[235:232] ^ 1);
  assign w884[20] = |(datain[231:228] ^ 10);
  assign w884[21] = |(datain[227:224] ^ 12);
  assign w884[22] = |(datain[223:220] ^ 3);
  assign w884[23] = |(datain[219:216] ^ 2);
  assign w884[24] = |(datain[215:212] ^ 12);
  assign w884[25] = |(datain[211:208] ^ 4);
  assign w884[26] = |(datain[207:204] ^ 14);
  assign w884[27] = |(datain[203:200] ^ 11);
  assign w884[28] = |(datain[199:196] ^ 0);
  assign w884[29] = |(datain[195:192] ^ 3);
  assign w884[30] = |(datain[191:188] ^ 9);
  assign w884[31] = |(datain[187:184] ^ 0);
  assign w884[32] = |(datain[183:180] ^ 15);
  assign w884[33] = |(datain[179:176] ^ 11);
  assign w884[34] = |(datain[175:172] ^ 13);
  assign w884[35] = |(datain[171:168] ^ 4);
  assign w884[36] = |(datain[167:164] ^ 10);
  assign w884[37] = |(datain[163:160] ^ 10);
  assign w884[38] = |(datain[159:156] ^ 14);
  assign w884[39] = |(datain[155:152] ^ 2);
  assign w884[40] = |(datain[151:148] ^ 15);
  assign w884[41] = |(datain[147:144] ^ 5);
  assign w884[42] = |(datain[143:140] ^ 14);
  assign w884[43] = |(datain[139:136] ^ 9);
  assign w884[44] = |(datain[135:132] ^ 10);
  assign w884[45] = |(datain[131:128] ^ 14);
  assign comp[884] = ~(|w884);
  wire [76-1:0] w885;
  assign w885[0] = |(datain[311:308] ^ 0);
  assign w885[1] = |(datain[307:304] ^ 4);
  assign w885[2] = |(datain[303:300] ^ 15);
  assign w885[3] = |(datain[299:296] ^ 10);
  assign w885[4] = |(datain[295:292] ^ 11);
  assign w885[5] = |(datain[291:288] ^ 14);
  assign w885[6] = |(datain[287:284] ^ 0);
  assign w885[7] = |(datain[283:280] ^ 0);
  assign w885[8] = |(datain[279:276] ^ 7);
  assign w885[9] = |(datain[275:272] ^ 12);
  assign w885[10] = |(datain[271:268] ^ 8);
  assign w885[11] = |(datain[267:264] ^ 14);
  assign w885[12] = |(datain[263:260] ^ 13);
  assign w885[13] = |(datain[259:256] ^ 7);
  assign w885[14] = |(datain[255:252] ^ 8);
  assign w885[15] = |(datain[251:248] ^ 11);
  assign w885[16] = |(datain[247:244] ^ 14);
  assign w885[17] = |(datain[243:240] ^ 6);
  assign w885[18] = |(datain[239:236] ^ 8);
  assign w885[19] = |(datain[235:232] ^ 14);
  assign w885[20] = |(datain[231:228] ^ 13);
  assign w885[21] = |(datain[227:224] ^ 15);
  assign w885[22] = |(datain[223:220] ^ 10);
  assign w885[23] = |(datain[219:216] ^ 1);
  assign w885[24] = |(datain[215:212] ^ 2);
  assign w885[25] = |(datain[211:208] ^ 2);
  assign w885[26] = |(datain[207:204] ^ 0);
  assign w885[27] = |(datain[203:200] ^ 0);
  assign w885[28] = |(datain[199:196] ^ 8);
  assign w885[29] = |(datain[195:192] ^ 0);
  assign w885[30] = |(datain[191:188] ^ 15);
  assign w885[31] = |(datain[187:184] ^ 12);
  assign w885[32] = |(datain[183:180] ^ 9);
  assign w885[33] = |(datain[179:176] ^ 15);
  assign w885[34] = |(datain[175:172] ^ 7);
  assign w885[35] = |(datain[171:168] ^ 4);
  assign w885[36] = |(datain[167:164] ^ 3);
  assign w885[37] = |(datain[163:160] ^ 11);
  assign w885[38] = |(datain[159:156] ^ 10);
  assign w885[39] = |(datain[155:152] ^ 3);
  assign w885[40] = |(datain[151:148] ^ 0);
  assign w885[41] = |(datain[147:144] ^ 6);
  assign w885[42] = |(datain[143:140] ^ 7);
  assign w885[43] = |(datain[139:136] ^ 12);
  assign w885[44] = |(datain[135:132] ^ 10);
  assign w885[45] = |(datain[131:128] ^ 1);
  assign w885[46] = |(datain[127:124] ^ 2);
  assign w885[47] = |(datain[123:120] ^ 0);
  assign w885[48] = |(datain[119:116] ^ 0);
  assign w885[49] = |(datain[115:112] ^ 0);
  assign w885[50] = |(datain[111:108] ^ 10);
  assign w885[51] = |(datain[107:104] ^ 3);
  assign w885[52] = |(datain[103:100] ^ 0);
  assign w885[53] = |(datain[99:96] ^ 4);
  assign w885[54] = |(datain[95:92] ^ 7);
  assign w885[55] = |(datain[91:88] ^ 12);
  assign w885[56] = |(datain[87:84] ^ 12);
  assign w885[57] = |(datain[83:80] ^ 4);
  assign w885[58] = |(datain[79:76] ^ 0);
  assign w885[59] = |(datain[75:72] ^ 6);
  assign w885[60] = |(datain[71:68] ^ 4);
  assign w885[61] = |(datain[67:64] ^ 12);
  assign w885[62] = |(datain[63:60] ^ 0);
  assign w885[63] = |(datain[59:56] ^ 0);
  assign w885[64] = |(datain[55:52] ^ 10);
  assign w885[65] = |(datain[51:48] ^ 3);
  assign w885[66] = |(datain[47:44] ^ 0);
  assign w885[67] = |(datain[43:40] ^ 8);
  assign w885[68] = |(datain[39:36] ^ 7);
  assign w885[69] = |(datain[35:32] ^ 12);
  assign w885[70] = |(datain[31:28] ^ 8);
  assign w885[71] = |(datain[27:24] ^ 12);
  assign w885[72] = |(datain[23:20] ^ 0);
  assign w885[73] = |(datain[19:16] ^ 6);
  assign w885[74] = |(datain[15:12] ^ 0);
  assign w885[75] = |(datain[11:8] ^ 10);
  assign comp[885] = ~(|w885);
  wire [46-1:0] w886;
  assign w886[0] = |(datain[311:308] ^ 2);
  assign w886[1] = |(datain[307:304] ^ 6);
  assign w886[2] = |(datain[303:300] ^ 0);
  assign w886[3] = |(datain[299:296] ^ 9);
  assign w886[4] = |(datain[295:292] ^ 0);
  assign w886[5] = |(datain[291:288] ^ 1);
  assign w886[6] = |(datain[287:284] ^ 11);
  assign w886[7] = |(datain[283:280] ^ 9);
  assign w886[8] = |(datain[279:276] ^ 12);
  assign w886[9] = |(datain[275:272] ^ 2);
  assign w886[10] = |(datain[271:268] ^ 0);
  assign w886[11] = |(datain[267:264] ^ 4);
  assign w886[12] = |(datain[263:260] ^ 11);
  assign w886[13] = |(datain[259:256] ^ 14);
  assign w886[14] = |(datain[255:252] ^ 0);
  assign w886[15] = |(datain[251:248] ^ 12);
  assign w886[16] = |(datain[247:244] ^ 0);
  assign w886[17] = |(datain[243:240] ^ 1);
  assign w886[18] = |(datain[239:236] ^ 8);
  assign w886[19] = |(datain[235:232] ^ 11);
  assign w886[20] = |(datain[231:228] ^ 15);
  assign w886[21] = |(datain[227:224] ^ 14);
  assign w886[22] = |(datain[223:220] ^ 15);
  assign w886[23] = |(datain[219:216] ^ 12);
  assign w886[24] = |(datain[215:212] ^ 10);
  assign w886[25] = |(datain[211:208] ^ 12);
  assign w886[26] = |(datain[207:204] ^ 3);
  assign w886[27] = |(datain[203:200] ^ 2);
  assign w886[28] = |(datain[199:196] ^ 12);
  assign w886[29] = |(datain[195:192] ^ 4);
  assign w886[30] = |(datain[191:188] ^ 10);
  assign w886[31] = |(datain[187:184] ^ 10);
  assign w886[32] = |(datain[183:180] ^ 14);
  assign w886[33] = |(datain[179:176] ^ 2);
  assign w886[34] = |(datain[175:172] ^ 15);
  assign w886[35] = |(datain[171:168] ^ 10);
  assign w886[36] = |(datain[167:164] ^ 12);
  assign w886[37] = |(datain[163:160] ^ 3);
  assign w886[38] = |(datain[159:156] ^ 0);
  assign w886[39] = |(datain[155:152] ^ 14);
  assign w886[40] = |(datain[151:148] ^ 0);
  assign w886[41] = |(datain[147:144] ^ 7);
  assign w886[42] = |(datain[143:140] ^ 0);
  assign w886[43] = |(datain[139:136] ^ 14);
  assign w886[44] = |(datain[135:132] ^ 1);
  assign w886[45] = |(datain[131:128] ^ 15);
  assign comp[886] = ~(|w886);
  wire [26-1:0] w887;
  assign w887[0] = |(datain[311:308] ^ 9);
  assign w887[1] = |(datain[307:304] ^ 0);
  assign w887[2] = |(datain[303:300] ^ 9);
  assign w887[3] = |(datain[299:296] ^ 0);
  assign w887[4] = |(datain[295:292] ^ 11);
  assign w887[5] = |(datain[291:288] ^ 9);
  assign w887[6] = |(datain[287:284] ^ 8);
  assign w887[7] = |(datain[283:280] ^ 0);
  assign w887[8] = |(datain[279:276] ^ 0);
  assign w887[9] = |(datain[275:272] ^ 0);
  assign w887[10] = |(datain[271:268] ^ 11);
  assign w887[11] = |(datain[267:264] ^ 14);
  assign w887[12] = |(datain[263:260] ^ 8);
  assign w887[13] = |(datain[259:256] ^ 0);
  assign w887[14] = |(datain[255:252] ^ 0);
  assign w887[15] = |(datain[251:248] ^ 0);
  assign w887[16] = |(datain[247:244] ^ 11);
  assign w887[17] = |(datain[243:240] ^ 15);
  assign w887[18] = |(datain[239:236] ^ 7);
  assign w887[19] = |(datain[235:232] ^ 15);
  assign w887[20] = |(datain[231:228] ^ 15);
  assign w887[21] = |(datain[227:224] ^ 15);
  assign w887[22] = |(datain[223:220] ^ 15);
  assign w887[23] = |(datain[219:216] ^ 3);
  assign w887[24] = |(datain[215:212] ^ 10);
  assign w887[25] = |(datain[211:208] ^ 4);
  assign comp[887] = ~(|w887);
  wire [32-1:0] w888;
  assign w888[0] = |(datain[311:308] ^ 11);
  assign w888[1] = |(datain[307:304] ^ 9);
  assign w888[2] = |(datain[303:300] ^ 8);
  assign w888[3] = |(datain[299:296] ^ 0);
  assign w888[4] = |(datain[295:292] ^ 0);
  assign w888[5] = |(datain[291:288] ^ 0);
  assign w888[6] = |(datain[287:284] ^ 11);
  assign w888[7] = |(datain[283:280] ^ 14);
  assign w888[8] = |(datain[279:276] ^ 7);
  assign w888[9] = |(datain[275:272] ^ 15);
  assign w888[10] = |(datain[271:268] ^ 15);
  assign w888[11] = |(datain[267:264] ^ 15);
  assign w888[12] = |(datain[263:260] ^ 11);
  assign w888[13] = |(datain[259:256] ^ 15);
  assign w888[14] = |(datain[255:252] ^ 8);
  assign w888[15] = |(datain[251:248] ^ 0);
  assign w888[16] = |(datain[247:244] ^ 0);
  assign w888[17] = |(datain[243:240] ^ 0);
  assign w888[18] = |(datain[239:236] ^ 15);
  assign w888[19] = |(datain[235:232] ^ 3);
  assign w888[20] = |(datain[231:228] ^ 10);
  assign w888[21] = |(datain[227:224] ^ 4);
  assign w888[22] = |(datain[223:220] ^ 11);
  assign w888[23] = |(datain[219:216] ^ 8);
  assign w888[24] = |(datain[215:212] ^ 15);
  assign w888[25] = |(datain[211:208] ^ 3);
  assign w888[26] = |(datain[207:204] ^ 10);
  assign w888[27] = |(datain[203:200] ^ 4);
  assign w888[28] = |(datain[199:196] ^ 10);
  assign w888[29] = |(datain[195:192] ^ 3);
  assign w888[30] = |(datain[191:188] ^ 15);
  assign w888[31] = |(datain[187:184] ^ 9);
  assign comp[888] = ~(|w888);
  wire [32-1:0] w889;
  assign w889[0] = |(datain[311:308] ^ 1);
  assign w889[1] = |(datain[307:304] ^ 14);
  assign w889[2] = |(datain[303:300] ^ 0);
  assign w889[3] = |(datain[299:296] ^ 14);
  assign w889[4] = |(datain[295:292] ^ 1);
  assign w889[5] = |(datain[291:288] ^ 15);
  assign w889[6] = |(datain[287:284] ^ 11);
  assign w889[7] = |(datain[283:280] ^ 4);
  assign w889[8] = |(datain[279:276] ^ 1);
  assign w889[9] = |(datain[275:272] ^ 9);
  assign w889[10] = |(datain[271:268] ^ 12);
  assign w889[11] = |(datain[267:264] ^ 13);
  assign w889[12] = |(datain[263:260] ^ 2);
  assign w889[13] = |(datain[259:256] ^ 1);
  assign w889[14] = |(datain[255:252] ^ 5);
  assign w889[15] = |(datain[251:248] ^ 0);
  assign w889[16] = |(datain[247:244] ^ 11);
  assign w889[17] = |(datain[243:240] ^ 2);
  assign w889[18] = |(datain[239:236] ^ 0);
  assign w889[19] = |(datain[235:232] ^ 2);
  assign w889[20] = |(datain[231:228] ^ 11);
  assign w889[21] = |(datain[227:224] ^ 4);
  assign w889[22] = |(datain[223:220] ^ 0);
  assign w889[23] = |(datain[219:216] ^ 14);
  assign w889[24] = |(datain[215:212] ^ 12);
  assign w889[25] = |(datain[211:208] ^ 13);
  assign w889[26] = |(datain[207:204] ^ 2);
  assign w889[27] = |(datain[203:200] ^ 1);
  assign w889[28] = |(datain[199:196] ^ 11);
  assign w889[29] = |(datain[195:192] ^ 4);
  assign w889[30] = |(datain[191:188] ^ 1);
  assign w889[31] = |(datain[187:184] ^ 10);
  assign comp[889] = ~(|w889);
  wire [42-1:0] w890;
  assign w890[0] = |(datain[311:308] ^ 0);
  assign w890[1] = |(datain[307:304] ^ 2);
  assign w890[2] = |(datain[303:300] ^ 11);
  assign w890[3] = |(datain[299:296] ^ 4);
  assign w890[4] = |(datain[295:292] ^ 0);
  assign w890[5] = |(datain[291:288] ^ 14);
  assign w890[6] = |(datain[287:284] ^ 12);
  assign w890[7] = |(datain[283:280] ^ 13);
  assign w890[8] = |(datain[279:276] ^ 2);
  assign w890[9] = |(datain[275:272] ^ 1);
  assign w890[10] = |(datain[271:268] ^ 11);
  assign w890[11] = |(datain[267:264] ^ 4);
  assign w890[12] = |(datain[263:260] ^ 1);
  assign w890[13] = |(datain[259:256] ^ 10);
  assign w890[14] = |(datain[255:252] ^ 11);
  assign w890[15] = |(datain[251:248] ^ 10);
  assign w890[16] = |(datain[247:244] ^ 0);
  assign w890[17] = |(datain[243:240] ^ 12);
  assign w890[18] = |(datain[239:236] ^ 0);
  assign w890[19] = |(datain[235:232] ^ 0);
  assign w890[20] = |(datain[231:228] ^ 0);
  assign w890[21] = |(datain[227:224] ^ 3);
  assign w890[22] = |(datain[223:220] ^ 13);
  assign w890[23] = |(datain[219:216] ^ 5);
  assign w890[24] = |(datain[215:212] ^ 12);
  assign w890[25] = |(datain[211:208] ^ 13);
  assign w890[26] = |(datain[207:204] ^ 2);
  assign w890[27] = |(datain[203:200] ^ 1);
  assign w890[28] = |(datain[199:196] ^ 11);
  assign w890[29] = |(datain[195:192] ^ 10);
  assign w890[30] = |(datain[191:188] ^ 0);
  assign w890[31] = |(datain[187:184] ^ 4);
  assign w890[32] = |(datain[183:180] ^ 0);
  assign w890[33] = |(datain[179:176] ^ 0);
  assign w890[34] = |(datain[175:172] ^ 0);
  assign w890[35] = |(datain[171:168] ^ 3);
  assign w890[36] = |(datain[167:164] ^ 13);
  assign w890[37] = |(datain[163:160] ^ 5);
  assign w890[38] = |(datain[159:156] ^ 11);
  assign w890[39] = |(datain[155:152] ^ 4);
  assign w890[40] = |(datain[151:148] ^ 4);
  assign w890[41] = |(datain[147:144] ^ 14);
  assign comp[890] = ~(|w890);
  wire [46-1:0] w891;
  assign w891[0] = |(datain[311:308] ^ 0);
  assign w891[1] = |(datain[307:304] ^ 1);
  assign w891[2] = |(datain[303:300] ^ 2);
  assign w891[3] = |(datain[299:296] ^ 5);
  assign w891[4] = |(datain[295:292] ^ 11);
  assign w891[5] = |(datain[291:288] ^ 10);
  assign w891[6] = |(datain[287:284] ^ 6);
  assign w891[7] = |(datain[283:280] ^ 0);
  assign w891[8] = |(datain[279:276] ^ 0);
  assign w891[9] = |(datain[275:272] ^ 1);
  assign w891[10] = |(datain[271:268] ^ 12);
  assign w891[11] = |(datain[267:264] ^ 13);
  assign w891[12] = |(datain[263:260] ^ 2);
  assign w891[13] = |(datain[259:256] ^ 1);
  assign w891[14] = |(datain[255:252] ^ 11);
  assign w891[15] = |(datain[251:248] ^ 0);
  assign w891[16] = |(datain[247:244] ^ 0);
  assign w891[17] = |(datain[243:240] ^ 3);
  assign w891[18] = |(datain[239:236] ^ 12);
  assign w891[19] = |(datain[235:232] ^ 13);
  assign w891[20] = |(datain[231:228] ^ 2);
  assign w891[21] = |(datain[227:224] ^ 1);
  assign w891[22] = |(datain[223:220] ^ 14);
  assign w891[23] = |(datain[219:216] ^ 11);
  assign w891[24] = |(datain[215:212] ^ 0);
  assign w891[25] = |(datain[211:208] ^ 3);
  assign w891[26] = |(datain[207:204] ^ 9);
  assign w891[27] = |(datain[203:200] ^ 0);
  assign w891[28] = |(datain[199:196] ^ 0);
  assign w891[29] = |(datain[195:192] ^ 0);
  assign w891[30] = |(datain[191:188] ^ 0);
  assign w891[31] = |(datain[187:184] ^ 0);
  assign w891[32] = |(datain[183:180] ^ 14);
  assign w891[33] = |(datain[179:176] ^ 8);
  assign w891[34] = |(datain[175:172] ^ 0);
  assign w891[35] = |(datain[171:168] ^ 3);
  assign w891[36] = |(datain[167:164] ^ 0);
  assign w891[37] = |(datain[163:160] ^ 0);
  assign w891[38] = |(datain[159:156] ^ 14);
  assign w891[39] = |(datain[155:152] ^ 11);
  assign w891[40] = |(datain[151:148] ^ 4);
  assign w891[41] = |(datain[147:144] ^ 7);
  assign w891[42] = |(datain[143:140] ^ 9);
  assign w891[43] = |(datain[139:136] ^ 0);
  assign w891[44] = |(datain[135:132] ^ 0);
  assign w891[45] = |(datain[131:128] ^ 14);
  assign comp[891] = ~(|w891);
  wire [48-1:0] w892;
  assign w892[0] = |(datain[311:308] ^ 3);
  assign w892[1] = |(datain[307:304] ^ 2);
  assign w892[2] = |(datain[303:300] ^ 12);
  assign w892[3] = |(datain[299:296] ^ 3);
  assign w892[4] = |(datain[295:292] ^ 10);
  assign w892[5] = |(datain[291:288] ^ 10);
  assign w892[6] = |(datain[287:284] ^ 14);
  assign w892[7] = |(datain[283:280] ^ 2);
  assign w892[8] = |(datain[279:276] ^ 15);
  assign w892[9] = |(datain[275:272] ^ 10);
  assign w892[10] = |(datain[271:268] ^ 2);
  assign w892[11] = |(datain[267:264] ^ 14);
  assign w892[12] = |(datain[263:260] ^ 8);
  assign w892[13] = |(datain[259:256] ^ 3);
  assign w892[14] = |(datain[255:252] ^ 3);
  assign w892[15] = |(datain[251:248] ^ 14);
  assign w892[16] = |(datain[247:244] ^ 0);
  assign w892[17] = |(datain[243:240] ^ 15);
  assign w892[18] = |(datain[239:236] ^ 0);
  assign w892[19] = |(datain[235:232] ^ 1);
  assign w892[20] = |(datain[231:228] ^ 0);
  assign w892[21] = |(datain[227:224] ^ 0);
  assign w892[22] = |(datain[223:220] ^ 7);
  assign w892[23] = |(datain[219:216] ^ 4);
  assign w892[24] = |(datain[215:212] ^ 2);
  assign w892[25] = |(datain[211:208] ^ 9);
  assign w892[26] = |(datain[207:204] ^ 11);
  assign w892[27] = |(datain[203:200] ^ 4);
  assign w892[28] = |(datain[199:196] ^ 4);
  assign w892[29] = |(datain[195:192] ^ 0);
  assign w892[30] = |(datain[191:188] ^ 2);
  assign w892[31] = |(datain[187:184] ^ 14);
  assign w892[32] = |(datain[183:180] ^ 8);
  assign w892[33] = |(datain[179:176] ^ 11);
  assign w892[34] = |(datain[175:172] ^ 1);
  assign w892[35] = |(datain[171:168] ^ 14);
  assign w892[36] = |(datain[167:164] ^ 0);
  assign w892[37] = |(datain[163:160] ^ 15);
  assign w892[38] = |(datain[159:156] ^ 0);
  assign w892[39] = |(datain[155:152] ^ 1);
  assign w892[40] = |(datain[151:148] ^ 2);
  assign w892[41] = |(datain[147:144] ^ 14);
  assign w892[42] = |(datain[143:140] ^ 15);
  assign w892[43] = |(datain[139:136] ^ 15);
  assign w892[44] = |(datain[135:132] ^ 3);
  assign w892[45] = |(datain[131:128] ^ 6);
  assign w892[46] = |(datain[127:124] ^ 0);
  assign w892[47] = |(datain[123:120] ^ 15);
  assign comp[892] = ~(|w892);
  wire [74-1:0] w893;
  assign w893[0] = |(datain[311:308] ^ 11);
  assign w893[1] = |(datain[307:304] ^ 9);
  assign w893[2] = |(datain[303:300] ^ 0);
  assign w893[3] = |(datain[299:296] ^ 3);
  assign w893[4] = |(datain[295:292] ^ 0);
  assign w893[5] = |(datain[291:288] ^ 0);
  assign w893[6] = |(datain[287:284] ^ 11);
  assign w893[7] = |(datain[283:280] ^ 10);
  assign w893[8] = |(datain[279:276] ^ 11);
  assign w893[9] = |(datain[275:272] ^ 6);
  assign w893[10] = |(datain[271:268] ^ 0);
  assign w893[11] = |(datain[267:264] ^ 2);
  assign w893[12] = |(datain[263:260] ^ 12);
  assign w893[13] = |(datain[259:256] ^ 13);
  assign w893[14] = |(datain[255:252] ^ 2);
  assign w893[15] = |(datain[251:248] ^ 1);
  assign w893[16] = |(datain[247:244] ^ 14);
  assign w893[17] = |(datain[243:240] ^ 8);
  assign w893[18] = |(datain[239:236] ^ 2);
  assign w893[19] = |(datain[235:232] ^ 6);
  assign w893[20] = |(datain[231:228] ^ 0);
  assign w893[21] = |(datain[227:224] ^ 0);
  assign w893[22] = |(datain[223:220] ^ 11);
  assign w893[23] = |(datain[219:216] ^ 4);
  assign w893[24] = |(datain[215:212] ^ 4);
  assign w893[25] = |(datain[211:208] ^ 0);
  assign w893[26] = |(datain[207:204] ^ 8);
  assign w893[27] = |(datain[203:200] ^ 11);
  assign w893[28] = |(datain[199:196] ^ 0);
  assign w893[29] = |(datain[195:192] ^ 14);
  assign w893[30] = |(datain[191:188] ^ 6);
  assign w893[31] = |(datain[187:184] ^ 2);
  assign w893[32] = |(datain[183:180] ^ 0);
  assign w893[33] = |(datain[179:176] ^ 1);
  assign w893[34] = |(datain[175:172] ^ 11);
  assign w893[35] = |(datain[171:168] ^ 10);
  assign w893[36] = |(datain[167:164] ^ 0);
  assign w893[37] = |(datain[163:160] ^ 0);
  assign w893[38] = |(datain[159:156] ^ 0);
  assign w893[39] = |(datain[155:152] ^ 1);
  assign w893[40] = |(datain[151:148] ^ 12);
  assign w893[41] = |(datain[147:144] ^ 13);
  assign w893[42] = |(datain[143:140] ^ 2);
  assign w893[43] = |(datain[139:136] ^ 1);
  assign w893[44] = |(datain[135:132] ^ 11);
  assign w893[45] = |(datain[131:128] ^ 4);
  assign w893[46] = |(datain[127:124] ^ 4);
  assign w893[47] = |(datain[123:120] ^ 0);
  assign w893[48] = |(datain[119:116] ^ 11);
  assign w893[49] = |(datain[115:112] ^ 9);
  assign w893[50] = |(datain[111:108] ^ 0);
  assign w893[51] = |(datain[107:104] ^ 3);
  assign w893[52] = |(datain[103:100] ^ 0);
  assign w893[53] = |(datain[99:96] ^ 0);
  assign w893[54] = |(datain[95:92] ^ 11);
  assign w893[55] = |(datain[91:88] ^ 10);
  assign w893[56] = |(datain[87:84] ^ 11);
  assign w893[57] = |(datain[83:80] ^ 9);
  assign w893[58] = |(datain[79:76] ^ 0);
  assign w893[59] = |(datain[75:72] ^ 2);
  assign w893[60] = |(datain[71:68] ^ 12);
  assign w893[61] = |(datain[67:64] ^ 13);
  assign w893[62] = |(datain[63:60] ^ 2);
  assign w893[63] = |(datain[59:56] ^ 1);
  assign w893[64] = |(datain[55:52] ^ 5);
  assign w893[65] = |(datain[51:48] ^ 9);
  assign w893[66] = |(datain[47:44] ^ 5);
  assign w893[67] = |(datain[43:40] ^ 10);
  assign w893[68] = |(datain[39:36] ^ 8);
  assign w893[69] = |(datain[35:32] ^ 0);
  assign w893[70] = |(datain[31:28] ^ 14);
  assign w893[71] = |(datain[27:24] ^ 1);
  assign w893[72] = |(datain[23:20] ^ 15);
  assign w893[73] = |(datain[19:16] ^ 0);
  assign comp[893] = ~(|w893);
  wire [32-1:0] w894;
  assign w894[0] = |(datain[311:308] ^ 3);
  assign w894[1] = |(datain[307:304] ^ 7);
  assign w894[2] = |(datain[303:300] ^ 5);
  assign w894[3] = |(datain[299:296] ^ 5);
  assign w894[4] = |(datain[295:292] ^ 7);
  assign w894[5] = |(datain[291:288] ^ 11);
  assign w894[6] = |(datain[287:284] ^ 7);
  assign w894[7] = |(datain[283:280] ^ 8);
  assign w894[8] = |(datain[279:276] ^ 7);
  assign w894[9] = |(datain[275:272] ^ 8);
  assign w894[10] = |(datain[271:268] ^ 7);
  assign w894[11] = |(datain[267:264] ^ 3);
  assign w894[12] = |(datain[263:260] ^ 6);
  assign w894[13] = |(datain[259:256] ^ 14);
  assign w894[14] = |(datain[255:252] ^ 3);
  assign w894[15] = |(datain[251:248] ^ 6);
  assign w894[16] = |(datain[247:244] ^ 3);
  assign w894[17] = |(datain[243:240] ^ 7);
  assign w894[18] = |(datain[239:236] ^ 5);
  assign w894[19] = |(datain[235:232] ^ 13);
  assign w894[20] = |(datain[231:228] ^ 6);
  assign w894[21] = |(datain[227:224] ^ 2);
  assign w894[22] = |(datain[223:220] ^ 7);
  assign w894[23] = |(datain[219:216] ^ 9);
  assign w894[24] = |(datain[215:212] ^ 3);
  assign w894[25] = |(datain[211:208] ^ 9);
  assign w894[26] = |(datain[207:204] ^ 3);
  assign w894[27] = |(datain[203:200] ^ 7);
  assign w894[28] = |(datain[199:196] ^ 2);
  assign w894[29] = |(datain[195:192] ^ 3);
  assign w894[30] = |(datain[191:188] ^ 3);
  assign w894[31] = |(datain[187:184] ^ 11);
  assign comp[894] = ~(|w894);
  wire [64-1:0] w895;
  assign w895[0] = |(datain[311:308] ^ 0);
  assign w895[1] = |(datain[307:304] ^ 2);
  assign w895[2] = |(datain[303:300] ^ 9);
  assign w895[3] = |(datain[299:296] ^ 0);
  assign w895[4] = |(datain[295:292] ^ 11);
  assign w895[5] = |(datain[291:288] ^ 11);
  assign w895[6] = |(datain[287:284] ^ 3);
  assign w895[7] = |(datain[283:280] ^ 11);
  assign w895[8] = |(datain[279:276] ^ 0);
  assign w895[9] = |(datain[275:272] ^ 1);
  assign w895[10] = |(datain[271:268] ^ 0);
  assign w895[11] = |(datain[267:264] ^ 3);
  assign w895[12] = |(datain[263:260] ^ 13);
  assign w895[13] = |(datain[259:256] ^ 14);
  assign w895[14] = |(datain[255:252] ^ 8);
  assign w895[15] = |(datain[251:248] ^ 10);
  assign w895[16] = |(datain[247:244] ^ 8);
  assign w895[17] = |(datain[243:240] ^ 4);
  assign w895[18] = |(datain[239:236] ^ 0);
  assign w895[19] = |(datain[235:232] ^ 12);
  assign w895[20] = |(datain[231:228] ^ 0);
  assign w895[21] = |(datain[227:224] ^ 1);
  assign w895[22] = |(datain[223:220] ^ 4);
  assign w895[23] = |(datain[219:216] ^ 15);
  assign w895[24] = |(datain[215:212] ^ 0);
  assign w895[25] = |(datain[211:208] ^ 4);
  assign w895[26] = |(datain[207:204] ^ 3);
  assign w895[27] = |(datain[203:200] ^ 0);
  assign w895[28] = |(datain[199:196] ^ 3);
  assign w895[29] = |(datain[195:192] ^ 0);
  assign w895[30] = |(datain[191:188] ^ 0);
  assign w895[31] = |(datain[187:184] ^ 1);
  assign w895[32] = |(datain[183:180] ^ 8);
  assign w895[33] = |(datain[179:176] ^ 3);
  assign w895[34] = |(datain[175:172] ^ 15);
  assign w895[35] = |(datain[171:168] ^ 15);
  assign w895[36] = |(datain[167:164] ^ 0);
  assign w895[37] = |(datain[163:160] ^ 0);
  assign w895[38] = |(datain[159:156] ^ 7);
  assign w895[39] = |(datain[155:152] ^ 5);
  assign w895[40] = |(datain[151:148] ^ 15);
  assign w895[41] = |(datain[147:144] ^ 6);
  assign w895[42] = |(datain[143:140] ^ 5);
  assign w895[43] = |(datain[139:136] ^ 11);
  assign w895[44] = |(datain[135:132] ^ 12);
  assign w895[45] = |(datain[131:128] ^ 3);
  assign w895[46] = |(datain[127:124] ^ 14);
  assign w895[47] = |(datain[123:120] ^ 8);
  assign w895[48] = |(datain[119:116] ^ 14);
  assign w895[49] = |(datain[115:112] ^ 3);
  assign w895[50] = |(datain[111:108] ^ 15);
  assign w895[51] = |(datain[107:104] ^ 15);
  assign w895[52] = |(datain[103:100] ^ 12);
  assign w895[53] = |(datain[99:96] ^ 13);
  assign w895[54] = |(datain[95:92] ^ 2);
  assign w895[55] = |(datain[91:88] ^ 1);
  assign w895[56] = |(datain[87:84] ^ 14);
  assign w895[57] = |(datain[83:80] ^ 8);
  assign w895[58] = |(datain[79:76] ^ 13);
  assign w895[59] = |(datain[75:72] ^ 14);
  assign w895[60] = |(datain[71:68] ^ 15);
  assign w895[61] = |(datain[67:64] ^ 15);
  assign w895[62] = |(datain[63:60] ^ 12);
  assign w895[63] = |(datain[59:56] ^ 3);
  assign comp[895] = ~(|w895);
  wire [74-1:0] w896;
  assign w896[0] = |(datain[311:308] ^ 3);
  assign w896[1] = |(datain[307:304] ^ 13);
  assign w896[2] = |(datain[303:300] ^ 4);
  assign w896[3] = |(datain[299:296] ^ 0);
  assign w896[4] = |(datain[295:292] ^ 3);
  assign w896[5] = |(datain[291:288] ^ 6);
  assign w896[6] = |(datain[287:284] ^ 9);
  assign w896[7] = |(datain[283:280] ^ 0);
  assign w896[8] = |(datain[279:276] ^ 0);
  assign w896[9] = |(datain[275:272] ^ 14);
  assign w896[10] = |(datain[271:268] ^ 1);
  assign w896[11] = |(datain[267:264] ^ 15);
  assign w896[12] = |(datain[263:260] ^ 8);
  assign w896[13] = |(datain[259:256] ^ 1);
  assign w896[14] = |(datain[255:252] ^ 7);
  assign w896[15] = |(datain[251:248] ^ 7);
  assign w896[16] = |(datain[247:244] ^ 2);
  assign w896[17] = |(datain[243:240] ^ 10);
  assign w896[18] = |(datain[239:236] ^ 4);
  assign w896[19] = |(datain[235:232] ^ 0);
  assign w896[20] = |(datain[231:228] ^ 3);
  assign w896[21] = |(datain[227:224] ^ 6);
  assign w896[22] = |(datain[223:220] ^ 9);
  assign w896[23] = |(datain[219:216] ^ 0);
  assign w896[24] = |(datain[215:212] ^ 8);
  assign w896[25] = |(datain[211:208] ^ 1);
  assign w896[26] = |(datain[207:204] ^ 7);
  assign w896[27] = |(datain[203:200] ^ 7);
  assign w896[28] = |(datain[199:196] ^ 2);
  assign w896[29] = |(datain[195:192] ^ 14);
  assign w896[30] = |(datain[191:188] ^ 4);
  assign w896[31] = |(datain[187:184] ^ 0);
  assign w896[32] = |(datain[183:180] ^ 3);
  assign w896[33] = |(datain[179:176] ^ 6);
  assign w896[34] = |(datain[175:172] ^ 9);
  assign w896[35] = |(datain[171:168] ^ 0);
  assign w896[36] = |(datain[167:164] ^ 8);
  assign w896[37] = |(datain[163:160] ^ 1);
  assign w896[38] = |(datain[159:156] ^ 7);
  assign w896[39] = |(datain[155:152] ^ 7);
  assign w896[40] = |(datain[151:148] ^ 3);
  assign w896[41] = |(datain[147:144] ^ 1);
  assign w896[42] = |(datain[143:140] ^ 4);
  assign w896[43] = |(datain[139:136] ^ 0);
  assign w896[44] = |(datain[135:132] ^ 3);
  assign w896[45] = |(datain[131:128] ^ 6);
  assign w896[46] = |(datain[127:124] ^ 9);
  assign w896[47] = |(datain[123:120] ^ 0);
  assign w896[48] = |(datain[119:116] ^ 8);
  assign w896[49] = |(datain[115:112] ^ 1);
  assign w896[50] = |(datain[111:108] ^ 7);
  assign w896[51] = |(datain[107:104] ^ 7);
  assign w896[52] = |(datain[103:100] ^ 3);
  assign w896[53] = |(datain[99:96] ^ 9);
  assign w896[54] = |(datain[95:92] ^ 4);
  assign w896[55] = |(datain[91:88] ^ 0);
  assign w896[56] = |(datain[87:84] ^ 3);
  assign w896[57] = |(datain[83:80] ^ 6);
  assign w896[58] = |(datain[79:76] ^ 9);
  assign w896[59] = |(datain[75:72] ^ 0);
  assign w896[60] = |(datain[71:68] ^ 8);
  assign w896[61] = |(datain[67:64] ^ 1);
  assign w896[62] = |(datain[63:60] ^ 7);
  assign w896[63] = |(datain[59:56] ^ 7);
  assign w896[64] = |(datain[55:52] ^ 3);
  assign w896[65] = |(datain[51:48] ^ 11);
  assign w896[66] = |(datain[47:44] ^ 4);
  assign w896[67] = |(datain[43:40] ^ 0);
  assign w896[68] = |(datain[39:36] ^ 3);
  assign w896[69] = |(datain[35:32] ^ 6);
  assign w896[70] = |(datain[31:28] ^ 9);
  assign w896[71] = |(datain[27:24] ^ 0);
  assign w896[72] = |(datain[23:20] ^ 15);
  assign w896[73] = |(datain[19:16] ^ 11);
  assign comp[896] = ~(|w896);
  wire [70-1:0] w897;
  assign w897[0] = |(datain[311:308] ^ 0);
  assign w897[1] = |(datain[307:304] ^ 3);
  assign w897[2] = |(datain[303:300] ^ 0);
  assign w897[3] = |(datain[299:296] ^ 0);
  assign w897[4] = |(datain[295:292] ^ 11);
  assign w897[5] = |(datain[291:288] ^ 9);
  assign w897[6] = |(datain[287:284] ^ 15);
  assign w897[7] = |(datain[283:280] ^ 15);
  assign w897[8] = |(datain[279:276] ^ 15);
  assign w897[9] = |(datain[275:272] ^ 15);
  assign w897[10] = |(datain[271:268] ^ 10);
  assign w897[11] = |(datain[267:264] ^ 12);
  assign w897[12] = |(datain[263:260] ^ 4);
  assign w897[13] = |(datain[259:256] ^ 9);
  assign w897[14] = |(datain[255:252] ^ 7);
  assign w897[15] = |(datain[251:248] ^ 5);
  assign w897[16] = |(datain[247:244] ^ 15);
  assign w897[17] = |(datain[243:240] ^ 13);
  assign w897[18] = |(datain[239:236] ^ 0);
  assign w897[19] = |(datain[235:232] ^ 14);
  assign w897[20] = |(datain[231:228] ^ 0);
  assign w897[21] = |(datain[227:224] ^ 14);
  assign w897[22] = |(datain[223:220] ^ 1);
  assign w897[23] = |(datain[219:216] ^ 15);
  assign w897[24] = |(datain[215:212] ^ 0);
  assign w897[25] = |(datain[211:208] ^ 7);
  assign w897[26] = |(datain[207:204] ^ 11);
  assign w897[27] = |(datain[203:200] ^ 14);
  assign w897[28] = |(datain[199:196] ^ 2);
  assign w897[29] = |(datain[195:192] ^ 10);
  assign w897[30] = |(datain[191:188] ^ 0);
  assign w897[31] = |(datain[187:184] ^ 0);
  assign w897[32] = |(datain[183:180] ^ 0);
  assign w897[33] = |(datain[179:176] ^ 3);
  assign w897[34] = |(datain[175:172] ^ 15);
  assign w897[35] = |(datain[171:168] ^ 5);
  assign w897[36] = |(datain[167:164] ^ 8);
  assign w897[37] = |(datain[163:160] ^ 11);
  assign w897[38] = |(datain[159:156] ^ 15);
  assign w897[39] = |(datain[155:152] ^ 14);
  assign w897[40] = |(datain[151:148] ^ 11);
  assign w897[41] = |(datain[147:144] ^ 9);
  assign w897[42] = |(datain[143:140] ^ 1);
  assign w897[43] = |(datain[139:136] ^ 3);
  assign w897[44] = |(datain[135:132] ^ 0);
  assign w897[45] = |(datain[131:128] ^ 4);
  assign w897[46] = |(datain[127:124] ^ 8);
  assign w897[47] = |(datain[123:120] ^ 10);
  assign w897[48] = |(datain[119:116] ^ 0);
  assign w897[49] = |(datain[115:112] ^ 4);
  assign w897[50] = |(datain[111:108] ^ 3);
  assign w897[51] = |(datain[107:104] ^ 4);
  assign w897[52] = |(datain[103:100] ^ 1);
  assign w897[53] = |(datain[99:96] ^ 2);
  assign w897[54] = |(datain[95:92] ^ 2);
  assign w897[55] = |(datain[91:88] ^ 6);
  assign w897[56] = |(datain[87:84] ^ 8);
  assign w897[57] = |(datain[83:80] ^ 8);
  assign w897[58] = |(datain[79:76] ^ 0);
  assign w897[59] = |(datain[75:72] ^ 5);
  assign w897[60] = |(datain[71:68] ^ 4);
  assign w897[61] = |(datain[67:64] ^ 6);
  assign w897[62] = |(datain[63:60] ^ 4);
  assign w897[63] = |(datain[59:56] ^ 7);
  assign w897[64] = |(datain[55:52] ^ 4);
  assign w897[65] = |(datain[51:48] ^ 9);
  assign w897[66] = |(datain[47:44] ^ 7);
  assign w897[67] = |(datain[43:40] ^ 5);
  assign w897[68] = |(datain[39:36] ^ 15);
  assign w897[69] = |(datain[35:32] ^ 4);
  assign comp[897] = ~(|w897);
  wire [76-1:0] w898;
  assign w898[0] = |(datain[311:308] ^ 3);
  assign w898[1] = |(datain[307:304] ^ 3);
  assign w898[2] = |(datain[303:300] ^ 12);
  assign w898[3] = |(datain[299:296] ^ 9);
  assign w898[4] = |(datain[295:292] ^ 3);
  assign w898[5] = |(datain[291:288] ^ 3);
  assign w898[6] = |(datain[287:284] ^ 13);
  assign w898[7] = |(datain[283:280] ^ 2);
  assign w898[8] = |(datain[279:276] ^ 14);
  assign w898[9] = |(datain[275:272] ^ 8);
  assign w898[10] = |(datain[271:268] ^ 2);
  assign w898[11] = |(datain[267:264] ^ 11);
  assign w898[12] = |(datain[263:260] ^ 0);
  assign w898[13] = |(datain[259:256] ^ 0);
  assign w898[14] = |(datain[255:252] ^ 12);
  assign w898[15] = |(datain[251:248] ^ 3);
  assign w898[16] = |(datain[247:244] ^ 5);
  assign w898[17] = |(datain[243:240] ^ 3);
  assign w898[18] = |(datain[239:236] ^ 11);
  assign w898[19] = |(datain[235:232] ^ 8);
  assign w898[20] = |(datain[231:228] ^ 11);
  assign w898[21] = |(datain[227:224] ^ 10);
  assign w898[22] = |(datain[223:220] ^ 1);
  assign w898[23] = |(datain[219:216] ^ 0);
  assign w898[24] = |(datain[215:212] ^ 3);
  assign w898[25] = |(datain[211:208] ^ 5);
  assign w898[26] = |(datain[207:204] ^ 9);
  assign w898[27] = |(datain[203:200] ^ 10);
  assign w898[28] = |(datain[199:196] ^ 0);
  assign w898[29] = |(datain[195:192] ^ 2);
  assign w898[30] = |(datain[191:188] ^ 12);
  assign w898[31] = |(datain[187:184] ^ 13);
  assign w898[32] = |(datain[183:180] ^ 2);
  assign w898[33] = |(datain[179:176] ^ 15);
  assign w898[34] = |(datain[175:172] ^ 7);
  assign w898[35] = |(datain[171:168] ^ 2);
  assign w898[36] = |(datain[167:164] ^ 1);
  assign w898[37] = |(datain[163:160] ^ 12);
  assign w898[38] = |(datain[159:156] ^ 2);
  assign w898[39] = |(datain[155:152] ^ 6);
  assign w898[40] = |(datain[151:148] ^ 8);
  assign w898[41] = |(datain[147:144] ^ 0);
  assign w898[42] = |(datain[143:140] ^ 3);
  assign w898[43] = |(datain[139:136] ^ 13);
  assign w898[44] = |(datain[135:132] ^ 15);
  assign w898[45] = |(datain[131:128] ^ 15);
  assign w898[46] = |(datain[127:124] ^ 7);
  assign w898[47] = |(datain[123:120] ^ 4);
  assign w898[48] = |(datain[119:116] ^ 1);
  assign w898[49] = |(datain[115:112] ^ 6);
  assign w898[50] = |(datain[111:108] ^ 3);
  assign w898[51] = |(datain[107:104] ^ 3);
  assign w898[52] = |(datain[103:100] ^ 13);
  assign w898[53] = |(datain[99:96] ^ 11);
  assign w898[54] = |(datain[95:92] ^ 2);
  assign w898[55] = |(datain[91:88] ^ 6);
  assign w898[56] = |(datain[87:84] ^ 8);
  assign w898[57] = |(datain[83:80] ^ 10);
  assign w898[58] = |(datain[79:76] ^ 1);
  assign w898[59] = |(datain[75:72] ^ 13);
  assign w898[60] = |(datain[71:68] ^ 11);
  assign w898[61] = |(datain[67:64] ^ 8);
  assign w898[62] = |(datain[63:60] ^ 8);
  assign w898[63] = |(datain[59:56] ^ 12);
  assign w898[64] = |(datain[55:52] ^ 1);
  assign w898[65] = |(datain[51:48] ^ 0);
  assign w898[66] = |(datain[47:44] ^ 3);
  assign w898[67] = |(datain[43:40] ^ 5);
  assign w898[68] = |(datain[39:36] ^ 9);
  assign w898[69] = |(datain[35:32] ^ 10);
  assign w898[70] = |(datain[31:28] ^ 0);
  assign w898[71] = |(datain[27:24] ^ 2);
  assign w898[72] = |(datain[23:20] ^ 12);
  assign w898[73] = |(datain[19:16] ^ 13);
  assign w898[74] = |(datain[15:12] ^ 2);
  assign w898[75] = |(datain[11:8] ^ 15);
  assign comp[898] = ~(|w898);
  wire [76-1:0] w899;
  assign w899[0] = |(datain[311:308] ^ 4);
  assign w899[1] = |(datain[307:304] ^ 13);
  assign w899[2] = |(datain[303:300] ^ 1);
  assign w899[3] = |(datain[299:296] ^ 2);
  assign w899[4] = |(datain[295:292] ^ 4);
  assign w899[5] = |(datain[291:288] ^ 3);
  assign w899[6] = |(datain[287:284] ^ 15);
  assign w899[7] = |(datain[283:280] ^ 14);
  assign w899[8] = |(datain[279:276] ^ 0);
  assign w899[9] = |(datain[275:272] ^ 6);
  assign w899[10] = |(datain[271:268] ^ 4);
  assign w899[11] = |(datain[267:264] ^ 15);
  assign w899[12] = |(datain[263:260] ^ 1);
  assign w899[13] = |(datain[259:256] ^ 2);
  assign w899[14] = |(datain[255:252] ^ 5);
  assign w899[15] = |(datain[251:248] ^ 0);
  assign w899[16] = |(datain[247:244] ^ 11);
  assign w899[17] = |(datain[243:240] ^ 4);
  assign w899[18] = |(datain[239:236] ^ 4);
  assign w899[19] = |(datain[235:232] ^ 0);
  assign w899[20] = |(datain[231:228] ^ 11);
  assign w899[21] = |(datain[227:224] ^ 9);
  assign w899[22] = |(datain[223:220] ^ 7);
  assign w899[23] = |(datain[219:216] ^ 13);
  assign w899[24] = |(datain[215:212] ^ 1);
  assign w899[25] = |(datain[211:208] ^ 2);
  assign w899[26] = |(datain[207:204] ^ 11);
  assign w899[27] = |(datain[203:200] ^ 10);
  assign w899[28] = |(datain[199:196] ^ 0);
  assign w899[29] = |(datain[195:192] ^ 0);
  assign w899[30] = |(datain[191:188] ^ 0);
  assign w899[31] = |(datain[187:184] ^ 0);
  assign w899[32] = |(datain[183:180] ^ 12);
  assign w899[33] = |(datain[179:176] ^ 13);
  assign w899[34] = |(datain[175:172] ^ 2);
  assign w899[35] = |(datain[171:168] ^ 1);
  assign w899[36] = |(datain[167:164] ^ 5);
  assign w899[37] = |(datain[163:160] ^ 8);
  assign w899[38] = |(datain[159:156] ^ 2);
  assign w899[39] = |(datain[155:152] ^ 13);
  assign w899[40] = |(datain[151:148] ^ 0);
  assign w899[41] = |(datain[147:144] ^ 3);
  assign w899[42] = |(datain[143:140] ^ 0);
  assign w899[43] = |(datain[139:136] ^ 0);
  assign w899[44] = |(datain[135:132] ^ 10);
  assign w899[45] = |(datain[131:128] ^ 3);
  assign w899[46] = |(datain[127:124] ^ 5);
  assign w899[47] = |(datain[123:120] ^ 9);
  assign w899[48] = |(datain[119:116] ^ 1);
  assign w899[49] = |(datain[115:112] ^ 2);
  assign w899[50] = |(datain[111:108] ^ 14);
  assign w899[51] = |(datain[107:104] ^ 8);
  assign w899[52] = |(datain[103:100] ^ 7);
  assign w899[53] = |(datain[99:96] ^ 2);
  assign w899[54] = |(datain[95:92] ^ 0);
  assign w899[55] = |(datain[91:88] ^ 4);
  assign w899[56] = |(datain[87:84] ^ 11);
  assign w899[57] = |(datain[83:80] ^ 4);
  assign w899[58] = |(datain[79:76] ^ 4);
  assign w899[59] = |(datain[75:72] ^ 0);
  assign w899[60] = |(datain[71:68] ^ 11);
  assign w899[61] = |(datain[67:64] ^ 9);
  assign w899[62] = |(datain[63:60] ^ 0);
  assign w899[63] = |(datain[59:56] ^ 5);
  assign w899[64] = |(datain[55:52] ^ 0);
  assign w899[65] = |(datain[51:48] ^ 0);
  assign w899[66] = |(datain[47:44] ^ 11);
  assign w899[67] = |(datain[43:40] ^ 10);
  assign w899[68] = |(datain[39:36] ^ 5);
  assign w899[69] = |(datain[35:32] ^ 8);
  assign w899[70] = |(datain[31:28] ^ 1);
  assign w899[71] = |(datain[27:24] ^ 2);
  assign w899[72] = |(datain[23:20] ^ 12);
  assign w899[73] = |(datain[19:16] ^ 13);
  assign w899[74] = |(datain[15:12] ^ 2);
  assign w899[75] = |(datain[11:8] ^ 1);
  assign comp[899] = ~(|w899);
  wire [76-1:0] w900;
  assign w900[0] = |(datain[311:308] ^ 0);
  assign w900[1] = |(datain[307:304] ^ 1);
  assign w900[2] = |(datain[303:300] ^ 11);
  assign w900[3] = |(datain[299:296] ^ 8);
  assign w900[4] = |(datain[295:292] ^ 0);
  assign w900[5] = |(datain[291:288] ^ 1);
  assign w900[6] = |(datain[287:284] ^ 0);
  assign w900[7] = |(datain[283:280] ^ 3);
  assign w900[8] = |(datain[279:276] ^ 11);
  assign w900[9] = |(datain[275:272] ^ 9);
  assign w900[10] = |(datain[271:268] ^ 0);
  assign w900[11] = |(datain[267:264] ^ 1);
  assign w900[12] = |(datain[263:260] ^ 0);
  assign w900[13] = |(datain[259:256] ^ 0);
  assign w900[14] = |(datain[255:252] ^ 12);
  assign w900[15] = |(datain[251:248] ^ 13);
  assign w900[16] = |(datain[247:244] ^ 1);
  assign w900[17] = |(datain[243:240] ^ 3);
  assign w900[18] = |(datain[239:236] ^ 5);
  assign w900[19] = |(datain[235:232] ^ 15);
  assign w900[20] = |(datain[231:228] ^ 5);
  assign w900[21] = |(datain[227:224] ^ 14);
  assign w900[22] = |(datain[223:220] ^ 5);
  assign w900[23] = |(datain[219:216] ^ 7);
  assign w900[24] = |(datain[215:212] ^ 11);
  assign w900[25] = |(datain[211:208] ^ 10);
  assign w900[26] = |(datain[207:204] ^ 6);
  assign w900[27] = |(datain[203:200] ^ 12);
  assign w900[28] = |(datain[199:196] ^ 0);
  assign w900[29] = |(datain[195:192] ^ 0);
  assign w900[30] = |(datain[191:188] ^ 0);
  assign w900[31] = |(datain[187:184] ^ 3);
  assign w900[32] = |(datain[183:180] ^ 13);
  assign w900[33] = |(datain[179:176] ^ 6);
  assign w900[34] = |(datain[175:172] ^ 11);
  assign w900[35] = |(datain[171:168] ^ 15);
  assign w900[36] = |(datain[167:164] ^ 8);
  assign w900[37] = |(datain[163:160] ^ 3);
  assign w900[38] = |(datain[159:156] ^ 0);
  assign w900[39] = |(datain[155:152] ^ 0);
  assign w900[40] = |(datain[151:148] ^ 0);
  assign w900[41] = |(datain[147:144] ^ 3);
  assign w900[42] = |(datain[143:140] ^ 15);
  assign w900[43] = |(datain[139:136] ^ 14);
  assign w900[44] = |(datain[135:132] ^ 11);
  assign w900[45] = |(datain[131:128] ^ 4);
  assign w900[46] = |(datain[127:124] ^ 5);
  assign w900[47] = |(datain[123:120] ^ 6);
  assign w900[48] = |(datain[119:116] ^ 12);
  assign w900[49] = |(datain[115:112] ^ 13);
  assign w900[50] = |(datain[111:108] ^ 2);
  assign w900[51] = |(datain[107:104] ^ 1);
  assign w900[52] = |(datain[103:100] ^ 11);
  assign w900[53] = |(datain[99:96] ^ 10);
  assign w900[54] = |(datain[95:92] ^ 7);
  assign w900[55] = |(datain[91:88] ^ 6);
  assign w900[56] = |(datain[87:84] ^ 0);
  assign w900[57] = |(datain[83:80] ^ 0);
  assign w900[58] = |(datain[79:76] ^ 0);
  assign w900[59] = |(datain[75:72] ^ 3);
  assign w900[60] = |(datain[71:68] ^ 13);
  assign w900[61] = |(datain[67:64] ^ 6);
  assign w900[62] = |(datain[63:60] ^ 11);
  assign w900[63] = |(datain[59:56] ^ 15);
  assign w900[64] = |(datain[55:52] ^ 9);
  assign w900[65] = |(datain[51:48] ^ 2);
  assign w900[66] = |(datain[47:44] ^ 0);
  assign w900[67] = |(datain[43:40] ^ 0);
  assign w900[68] = |(datain[39:36] ^ 0);
  assign w900[69] = |(datain[35:32] ^ 3);
  assign w900[70] = |(datain[31:28] ^ 15);
  assign w900[71] = |(datain[27:24] ^ 14);
  assign w900[72] = |(datain[23:20] ^ 11);
  assign w900[73] = |(datain[19:16] ^ 4);
  assign w900[74] = |(datain[15:12] ^ 5);
  assign w900[75] = |(datain[11:8] ^ 6);
  assign comp[900] = ~(|w900);
  wire [74-1:0] w901;
  assign w901[0] = |(datain[311:308] ^ 12);
  assign w901[1] = |(datain[307:304] ^ 13);
  assign w901[2] = |(datain[303:300] ^ 1);
  assign w901[3] = |(datain[299:296] ^ 3);
  assign w901[4] = |(datain[295:292] ^ 10);
  assign w901[5] = |(datain[291:288] ^ 1);
  assign w901[6] = |(datain[287:284] ^ 11);
  assign w901[7] = |(datain[283:280] ^ 12);
  assign w901[8] = |(datain[279:276] ^ 0);
  assign w901[9] = |(datain[275:272] ^ 3);
  assign w901[10] = |(datain[271:268] ^ 3);
  assign w901[11] = |(datain[267:264] ^ 13);
  assign w901[12] = |(datain[263:260] ^ 5);
  assign w901[13] = |(datain[259:256] ^ 0);
  assign w901[14] = |(datain[255:252] ^ 6);
  assign w901[15] = |(datain[251:248] ^ 8);
  assign w901[16] = |(datain[247:244] ^ 7);
  assign w901[17] = |(datain[243:240] ^ 4);
  assign w901[18] = |(datain[239:236] ^ 1);
  assign w901[19] = |(datain[235:232] ^ 10);
  assign w901[20] = |(datain[231:228] ^ 11);
  assign w901[21] = |(datain[227:224] ^ 15);
  assign w901[22] = |(datain[223:220] ^ 11);
  assign w901[23] = |(datain[219:216] ^ 12);
  assign w901[24] = |(datain[215:212] ^ 0);
  assign w901[25] = |(datain[211:208] ^ 3);
  assign w901[26] = |(datain[207:204] ^ 11);
  assign w901[27] = |(datain[203:200] ^ 8);
  assign w901[28] = |(datain[199:196] ^ 5);
  assign w901[29] = |(datain[195:192] ^ 4);
  assign w901[30] = |(datain[191:188] ^ 0);
  assign w901[31] = |(datain[187:184] ^ 0);
  assign w901[32] = |(datain[183:180] ^ 0);
  assign w901[33] = |(datain[179:176] ^ 3);
  assign w901[34] = |(datain[175:172] ^ 12);
  assign w901[35] = |(datain[171:168] ^ 6);
  assign w901[36] = |(datain[167:164] ^ 5);
  assign w901[37] = |(datain[163:160] ^ 0);
  assign w901[38] = |(datain[159:156] ^ 5);
  assign w901[39] = |(datain[155:152] ^ 14);
  assign w901[40] = |(datain[151:148] ^ 11);
  assign w901[41] = |(datain[147:144] ^ 9);
  assign w901[42] = |(datain[143:140] ^ 1);
  assign w901[43] = |(datain[139:136] ^ 7);
  assign w901[44] = |(datain[135:132] ^ 0);
  assign w901[45] = |(datain[131:128] ^ 0);
  assign w901[46] = |(datain[127:124] ^ 15);
  assign w901[47] = |(datain[123:120] ^ 3);
  assign w901[48] = |(datain[119:116] ^ 10);
  assign w901[49] = |(datain[115:112] ^ 4);
  assign w901[50] = |(datain[111:108] ^ 11);
  assign w901[51] = |(datain[107:104] ^ 10);
  assign w901[52] = |(datain[103:100] ^ 8);
  assign w901[53] = |(datain[99:96] ^ 0);
  assign w901[54] = |(datain[95:92] ^ 0);
  assign w901[55] = |(datain[91:88] ^ 0);
  assign w901[56] = |(datain[87:84] ^ 11);
  assign w901[57] = |(datain[83:80] ^ 8);
  assign w901[58] = |(datain[79:76] ^ 0);
  assign w901[59] = |(datain[75:72] ^ 1);
  assign w901[60] = |(datain[71:68] ^ 0);
  assign w901[61] = |(datain[67:64] ^ 3);
  assign w901[62] = |(datain[63:60] ^ 11);
  assign w901[63] = |(datain[59:56] ^ 9);
  assign w901[64] = |(datain[55:52] ^ 0);
  assign w901[65] = |(datain[51:48] ^ 1);
  assign w901[66] = |(datain[47:44] ^ 0);
  assign w901[67] = |(datain[43:40] ^ 0);
  assign w901[68] = |(datain[39:36] ^ 12);
  assign w901[69] = |(datain[35:32] ^ 13);
  assign w901[70] = |(datain[31:28] ^ 1);
  assign w901[71] = |(datain[27:24] ^ 3);
  assign w901[72] = |(datain[23:20] ^ 5);
  assign w901[73] = |(datain[19:16] ^ 15);
  assign comp[901] = ~(|w901);
  wire [42-1:0] w902;
  assign w902[0] = |(datain[311:308] ^ 8);
  assign w902[1] = |(datain[307:304] ^ 3);
  assign w902[2] = |(datain[303:300] ^ 12);
  assign w902[3] = |(datain[299:296] ^ 6);
  assign w902[4] = |(datain[295:292] ^ 1);
  assign w902[5] = |(datain[291:288] ^ 9);
  assign w902[6] = |(datain[287:284] ^ 11);
  assign w902[7] = |(datain[283:280] ^ 15);
  assign w902[8] = |(datain[279:276] ^ 0);
  assign w902[9] = |(datain[275:272] ^ 0);
  assign w902[10] = |(datain[271:268] ^ 0);
  assign w902[11] = |(datain[267:264] ^ 1);
  assign w902[12] = |(datain[263:260] ^ 11);
  assign w902[13] = |(datain[259:256] ^ 9);
  assign w902[14] = |(datain[255:252] ^ 0);
  assign w902[15] = |(datain[251:248] ^ 3);
  assign w902[16] = |(datain[247:244] ^ 0);
  assign w902[17] = |(datain[243:240] ^ 0);
  assign w902[18] = |(datain[239:236] ^ 15);
  assign w902[19] = |(datain[235:232] ^ 3);
  assign w902[20] = |(datain[231:228] ^ 10);
  assign w902[21] = |(datain[227:224] ^ 4);
  assign w902[22] = |(datain[223:220] ^ 8);
  assign w902[23] = |(datain[219:216] ^ 11);
  assign w902[24] = |(datain[215:212] ^ 15);
  assign w902[25] = |(datain[211:208] ^ 2);
  assign w902[26] = |(datain[207:204] ^ 11);
  assign w902[27] = |(datain[203:200] ^ 8);
  assign w902[28] = |(datain[199:196] ^ 2);
  assign w902[29] = |(datain[195:192] ^ 4);
  assign w902[30] = |(datain[191:188] ^ 3);
  assign w902[31] = |(datain[187:184] ^ 5);
  assign w902[32] = |(datain[183:180] ^ 12);
  assign w902[33] = |(datain[179:176] ^ 13);
  assign w902[34] = |(datain[175:172] ^ 2);
  assign w902[35] = |(datain[171:168] ^ 1);
  assign w902[36] = |(datain[167:164] ^ 0);
  assign w902[37] = |(datain[163:160] ^ 6);
  assign w902[38] = |(datain[159:156] ^ 5);
  assign w902[39] = |(datain[155:152] ^ 3);
  assign w902[40] = |(datain[151:148] ^ 11);
  assign w902[41] = |(datain[147:144] ^ 8);
  assign comp[902] = ~(|w902);
  wire [44-1:0] w903;
  assign w903[0] = |(datain[311:308] ^ 0);
  assign w903[1] = |(datain[307:304] ^ 14);
  assign w903[2] = |(datain[303:300] ^ 15);
  assign w903[3] = |(datain[299:296] ^ 14);
  assign w903[4] = |(datain[295:292] ^ 0);
  assign w903[5] = |(datain[291:288] ^ 1);
  assign w903[6] = |(datain[287:284] ^ 2);
  assign w903[7] = |(datain[283:280] ^ 6);
  assign w903[8] = |(datain[279:276] ^ 8);
  assign w903[9] = |(datain[275:272] ^ 11);
  assign w903[10] = |(datain[271:268] ^ 1);
  assign w903[11] = |(datain[267:264] ^ 14);
  assign w903[12] = |(datain[263:260] ^ 15);
  assign w903[13] = |(datain[259:256] ^ 12);
  assign w903[14] = |(datain[255:252] ^ 0);
  assign w903[15] = |(datain[251:248] ^ 1);
  assign w903[16] = |(datain[247:244] ^ 8);
  assign w903[17] = |(datain[243:240] ^ 3);
  assign w903[18] = |(datain[239:236] ^ 12);
  assign w903[19] = |(datain[235:232] ^ 1);
  assign w903[20] = |(datain[231:228] ^ 0);
  assign w903[21] = |(datain[227:224] ^ 1);
  assign w903[22] = |(datain[223:220] ^ 15);
  assign w903[23] = |(datain[219:216] ^ 10);
  assign w903[24] = |(datain[215:212] ^ 2);
  assign w903[25] = |(datain[211:208] ^ 6);
  assign w903[26] = |(datain[207:204] ^ 2);
  assign w903[27] = |(datain[203:200] ^ 11);
  assign w903[28] = |(datain[199:196] ^ 1);
  assign w903[29] = |(datain[195:192] ^ 14);
  assign w903[30] = |(datain[191:188] ^ 6);
  assign w903[31] = |(datain[187:184] ^ 12);
  assign w903[32] = |(datain[183:180] ^ 0);
  assign w903[33] = |(datain[179:176] ^ 4);
  assign w903[34] = |(datain[175:172] ^ 2);
  assign w903[35] = |(datain[171:168] ^ 6);
  assign w903[36] = |(datain[167:164] ^ 1);
  assign w903[37] = |(datain[163:160] ^ 11);
  assign w903[38] = |(datain[159:156] ^ 0);
  assign w903[39] = |(datain[155:152] ^ 14);
  assign w903[40] = |(datain[151:148] ^ 6);
  assign w903[41] = |(datain[147:144] ^ 14);
  assign w903[42] = |(datain[143:140] ^ 0);
  assign w903[43] = |(datain[139:136] ^ 4);
  assign comp[903] = ~(|w903);
  wire [28-1:0] w904;
  assign w904[0] = |(datain[311:308] ^ 0);
  assign w904[1] = |(datain[307:304] ^ 2);
  assign w904[2] = |(datain[303:300] ^ 4);
  assign w904[3] = |(datain[299:296] ^ 2);
  assign w904[4] = |(datain[295:292] ^ 12);
  assign w904[5] = |(datain[291:288] ^ 13);
  assign w904[6] = |(datain[287:284] ^ 2);
  assign w904[7] = |(datain[283:280] ^ 1);
  assign w904[8] = |(datain[279:276] ^ 11);
  assign w904[9] = |(datain[275:272] ^ 9);
  assign w904[10] = |(datain[271:268] ^ 11);
  assign w904[11] = |(datain[267:264] ^ 10);
  assign w904[12] = |(datain[263:260] ^ 0);
  assign w904[13] = |(datain[259:256] ^ 2);
  assign w904[14] = |(datain[255:252] ^ 11);
  assign w904[15] = |(datain[251:248] ^ 4);
  assign w904[16] = |(datain[247:244] ^ 4);
  assign w904[17] = |(datain[243:240] ^ 0);
  assign w904[18] = |(datain[239:236] ^ 11);
  assign w904[19] = |(datain[235:232] ^ 10);
  assign w904[20] = |(datain[231:228] ^ 12);
  assign w904[21] = |(datain[227:224] ^ 0);
  assign w904[22] = |(datain[223:220] ^ 0);
  assign w904[23] = |(datain[219:216] ^ 0);
  assign w904[24] = |(datain[215:212] ^ 12);
  assign w904[25] = |(datain[211:208] ^ 13);
  assign w904[26] = |(datain[207:204] ^ 2);
  assign w904[27] = |(datain[203:200] ^ 1);
  assign comp[904] = ~(|w904);
  wire [46-1:0] w905;
  assign w905[0] = |(datain[311:308] ^ 0);
  assign w905[1] = |(datain[307:304] ^ 6);
  assign w905[2] = |(datain[303:300] ^ 8);
  assign w905[3] = |(datain[299:296] ^ 0);
  assign w905[4] = |(datain[295:292] ^ 15);
  assign w905[5] = |(datain[291:288] ^ 12);
  assign w905[6] = |(datain[287:284] ^ 15);
  assign w905[7] = |(datain[283:280] ^ 14);
  assign w905[8] = |(datain[279:276] ^ 7);
  assign w905[9] = |(datain[275:272] ^ 5);
  assign w905[10] = |(datain[271:268] ^ 0);
  assign w905[11] = |(datain[267:264] ^ 15);
  assign w905[12] = |(datain[263:260] ^ 8);
  assign w905[13] = |(datain[259:256] ^ 1);
  assign w905[14] = |(datain[255:252] ^ 15);
  assign w905[15] = |(datain[251:248] ^ 11);
  assign w905[16] = |(datain[247:244] ^ 5);
  assign w905[17] = |(datain[243:240] ^ 2);
  assign w905[18] = |(datain[239:236] ^ 5);
  assign w905[19] = |(datain[235:232] ^ 3);
  assign w905[20] = |(datain[231:228] ^ 7);
  assign w905[21] = |(datain[227:224] ^ 4);
  assign w905[22] = |(datain[223:220] ^ 0);
  assign w905[23] = |(datain[219:216] ^ 3);
  assign w905[24] = |(datain[215:212] ^ 14);
  assign w905[25] = |(datain[211:208] ^ 9);
  assign w905[26] = |(datain[207:204] ^ 2);
  assign w905[27] = |(datain[203:200] ^ 8);
  assign w905[28] = |(datain[199:196] ^ 0);
  assign w905[29] = |(datain[195:192] ^ 1);
  assign w905[30] = |(datain[191:188] ^ 0);
  assign w905[31] = |(datain[187:184] ^ 7);
  assign w905[32] = |(datain[183:180] ^ 1);
  assign w905[33] = |(datain[179:176] ^ 15);
  assign w905[34] = |(datain[175:172] ^ 6);
  assign w905[35] = |(datain[171:168] ^ 1);
  assign w905[36] = |(datain[167:164] ^ 8);
  assign w905[37] = |(datain[163:160] ^ 11);
  assign w905[38] = |(datain[159:156] ^ 12);
  assign w905[39] = |(datain[155:152] ^ 3);
  assign w905[40] = |(datain[151:148] ^ 12);
  assign w905[41] = |(datain[147:144] ^ 15);
  assign w905[42] = |(datain[143:140] ^ 8);
  assign w905[43] = |(datain[139:136] ^ 0);
  assign w905[44] = |(datain[135:132] ^ 15);
  assign w905[45] = |(datain[131:128] ^ 12);
  assign comp[905] = ~(|w905);
  wire [76-1:0] w906;
  assign w906[0] = |(datain[311:308] ^ 2);
  assign w906[1] = |(datain[307:304] ^ 5);
  assign w906[2] = |(datain[303:300] ^ 11);
  assign w906[3] = |(datain[299:296] ^ 10);
  assign w906[4] = |(datain[295:292] ^ 11);
  assign w906[5] = |(datain[291:288] ^ 7);
  assign w906[6] = |(datain[287:284] ^ 0);
  assign w906[7] = |(datain[283:280] ^ 1);
  assign w906[8] = |(datain[279:276] ^ 9);
  assign w906[9] = |(datain[275:272] ^ 12);
  assign w906[10] = |(datain[271:268] ^ 15);
  assign w906[11] = |(datain[267:264] ^ 15);
  assign w906[12] = |(datain[263:260] ^ 1);
  assign w906[13] = |(datain[259:256] ^ 14);
  assign w906[14] = |(datain[255:252] ^ 3);
  assign w906[15] = |(datain[251:248] ^ 3);
  assign w906[16] = |(datain[247:244] ^ 0);
  assign w906[17] = |(datain[243:240] ^ 0);
  assign w906[18] = |(datain[239:236] ^ 11);
  assign w906[19] = |(datain[235:232] ^ 4);
  assign w906[20] = |(datain[231:228] ^ 4);
  assign w906[21] = |(datain[227:224] ^ 0);
  assign w906[22] = |(datain[223:220] ^ 11);
  assign w906[23] = |(datain[219:216] ^ 9);
  assign w906[24] = |(datain[215:212] ^ 2);
  assign w906[25] = |(datain[211:208] ^ 14);
  assign w906[26] = |(datain[207:204] ^ 0);
  assign w906[27] = |(datain[203:200] ^ 3);
  assign w906[28] = |(datain[199:196] ^ 3);
  assign w906[29] = |(datain[195:192] ^ 3);
  assign w906[30] = |(datain[191:188] ^ 13);
  assign w906[31] = |(datain[187:184] ^ 2);
  assign w906[32] = |(datain[183:180] ^ 9);
  assign w906[33] = |(datain[179:176] ^ 12);
  assign w906[34] = |(datain[175:172] ^ 15);
  assign w906[35] = |(datain[171:168] ^ 15);
  assign w906[36] = |(datain[167:164] ^ 1);
  assign w906[37] = |(datain[163:160] ^ 14);
  assign w906[38] = |(datain[159:156] ^ 3);
  assign w906[39] = |(datain[155:152] ^ 3);
  assign w906[40] = |(datain[151:148] ^ 0);
  assign w906[41] = |(datain[147:144] ^ 0);
  assign w906[42] = |(datain[143:140] ^ 11);
  assign w906[43] = |(datain[139:136] ^ 8);
  assign w906[44] = |(datain[135:132] ^ 0);
  assign w906[45] = |(datain[131:128] ^ 2);
  assign w906[46] = |(datain[127:124] ^ 4);
  assign w906[47] = |(datain[123:120] ^ 2);
  assign w906[48] = |(datain[119:116] ^ 8);
  assign w906[49] = |(datain[115:112] ^ 11);
  assign w906[50] = |(datain[111:108] ^ 12);
  assign w906[51] = |(datain[107:104] ^ 10);
  assign w906[52] = |(datain[103:100] ^ 9);
  assign w906[53] = |(datain[99:96] ^ 12);
  assign w906[54] = |(datain[95:92] ^ 15);
  assign w906[55] = |(datain[91:88] ^ 15);
  assign w906[56] = |(datain[87:84] ^ 1);
  assign w906[57] = |(datain[83:80] ^ 14);
  assign w906[58] = |(datain[79:76] ^ 3);
  assign w906[59] = |(datain[75:72] ^ 3);
  assign w906[60] = |(datain[71:68] ^ 0);
  assign w906[61] = |(datain[67:64] ^ 0);
  assign w906[62] = |(datain[63:60] ^ 8);
  assign w906[63] = |(datain[59:56] ^ 10);
  assign w906[64] = |(datain[55:52] ^ 15);
  assign w906[65] = |(datain[51:48] ^ 2);
  assign w906[66] = |(datain[47:44] ^ 8);
  assign w906[67] = |(datain[43:40] ^ 10);
  assign w906[68] = |(datain[39:36] ^ 13);
  assign w906[69] = |(datain[35:32] ^ 4);
  assign w906[70] = |(datain[31:28] ^ 13);
  assign w906[71] = |(datain[27:24] ^ 1);
  assign w906[72] = |(datain[23:20] ^ 14);
  assign w906[73] = |(datain[19:16] ^ 10);
  assign w906[74] = |(datain[15:12] ^ 10);
  assign w906[75] = |(datain[11:8] ^ 9);
  assign comp[906] = ~(|w906);
  wire [74-1:0] w907;
  assign w907[0] = |(datain[311:308] ^ 8);
  assign w907[1] = |(datain[307:304] ^ 11);
  assign w907[2] = |(datain[303:300] ^ 15);
  assign w907[3] = |(datain[299:296] ^ 5);
  assign w907[4] = |(datain[295:292] ^ 10);
  assign w907[5] = |(datain[291:288] ^ 4);
  assign w907[6] = |(datain[287:284] ^ 10);
  assign w907[7] = |(datain[283:280] ^ 4);
  assign w907[8] = |(datain[279:276] ^ 10);
  assign w907[9] = |(datain[275:272] ^ 4);
  assign w907[10] = |(datain[271:268] ^ 11);
  assign w907[11] = |(datain[267:264] ^ 8);
  assign w907[12] = |(datain[263:260] ^ 10);
  assign w907[13] = |(datain[259:256] ^ 11);
  assign w907[14] = |(datain[255:252] ^ 4);
  assign w907[15] = |(datain[251:248] ^ 11);
  assign w907[16] = |(datain[247:244] ^ 12);
  assign w907[17] = |(datain[243:240] ^ 13);
  assign w907[18] = |(datain[239:236] ^ 2);
  assign w907[19] = |(datain[235:232] ^ 1);
  assign w907[20] = |(datain[231:228] ^ 3);
  assign w907[21] = |(datain[227:224] ^ 13);
  assign w907[22] = |(datain[223:220] ^ 11);
  assign w907[23] = |(datain[219:216] ^ 0);
  assign w907[24] = |(datain[215:212] ^ 11);
  assign w907[25] = |(datain[211:208] ^ 0);
  assign w907[26] = |(datain[207:204] ^ 7);
  assign w907[27] = |(datain[203:200] ^ 5);
  assign w907[28] = |(datain[199:196] ^ 1);
  assign w907[29] = |(datain[195:192] ^ 7);
  assign w907[30] = |(datain[191:188] ^ 0);
  assign w907[31] = |(datain[187:184] ^ 14);
  assign w907[32] = |(datain[183:180] ^ 1);
  assign w907[33] = |(datain[179:176] ^ 15);
  assign w907[34] = |(datain[175:172] ^ 0);
  assign w907[35] = |(datain[171:168] ^ 14);
  assign w907[36] = |(datain[167:164] ^ 0);
  assign w907[37] = |(datain[163:160] ^ 7);
  assign w907[38] = |(datain[159:156] ^ 3);
  assign w907[39] = |(datain[155:152] ^ 3);
  assign w907[40] = |(datain[151:148] ^ 12);
  assign w907[41] = |(datain[147:144] ^ 0);
  assign w907[42] = |(datain[143:140] ^ 3);
  assign w907[43] = |(datain[139:136] ^ 3);
  assign w907[44] = |(datain[135:132] ^ 13);
  assign w907[45] = |(datain[131:128] ^ 11);
  assign w907[46] = |(datain[127:124] ^ 3);
  assign w907[47] = |(datain[123:120] ^ 3);
  assign w907[48] = |(datain[119:116] ^ 12);
  assign w907[49] = |(datain[115:112] ^ 9);
  assign w907[50] = |(datain[111:108] ^ 3);
  assign w907[51] = |(datain[107:104] ^ 3);
  assign w907[52] = |(datain[103:100] ^ 13);
  assign w907[53] = |(datain[99:96] ^ 2);
  assign w907[54] = |(datain[95:92] ^ 3);
  assign w907[55] = |(datain[91:88] ^ 3);
  assign w907[56] = |(datain[87:84] ^ 14);
  assign w907[57] = |(datain[83:80] ^ 13);
  assign w907[58] = |(datain[79:76] ^ 3);
  assign w907[59] = |(datain[75:72] ^ 3);
  assign w907[60] = |(datain[71:68] ^ 15);
  assign w907[61] = |(datain[67:64] ^ 15);
  assign w907[62] = |(datain[63:60] ^ 11);
  assign w907[63] = |(datain[59:56] ^ 14);
  assign w907[64] = |(datain[55:52] ^ 0);
  assign w907[65] = |(datain[51:48] ^ 0);
  assign w907[66] = |(datain[47:44] ^ 0);
  assign w907[67] = |(datain[43:40] ^ 1);
  assign w907[68] = |(datain[39:36] ^ 5);
  assign w907[69] = |(datain[35:32] ^ 6);
  assign w907[70] = |(datain[31:28] ^ 3);
  assign w907[71] = |(datain[27:24] ^ 3);
  assign w907[72] = |(datain[23:20] ^ 15);
  assign w907[73] = |(datain[19:16] ^ 6);
  assign comp[907] = ~(|w907);
  wire [42-1:0] w908;
  assign w908[0] = |(datain[311:308] ^ 0);
  assign w908[1] = |(datain[307:304] ^ 7);
  assign w908[2] = |(datain[303:300] ^ 7);
  assign w908[3] = |(datain[299:296] ^ 2);
  assign w908[4] = |(datain[295:292] ^ 0);
  assign w908[5] = |(datain[291:288] ^ 6);
  assign w908[6] = |(datain[287:284] ^ 8);
  assign w908[7] = |(datain[283:280] ^ 0);
  assign w908[8] = |(datain[279:276] ^ 15);
  assign w908[9] = |(datain[275:272] ^ 14);
  assign w908[10] = |(datain[271:268] ^ 0);
  assign w908[11] = |(datain[267:264] ^ 1);
  assign w908[12] = |(datain[263:260] ^ 7);
  assign w908[13] = |(datain[259:256] ^ 5);
  assign w908[14] = |(datain[255:252] ^ 0);
  assign w908[15] = |(datain[251:248] ^ 1);
  assign w908[16] = |(datain[247:244] ^ 4);
  assign w908[17] = |(datain[243:240] ^ 5);
  assign w908[18] = |(datain[239:236] ^ 11);
  assign w908[19] = |(datain[235:232] ^ 2);
  assign w908[20] = |(datain[231:228] ^ 0);
  assign w908[21] = |(datain[227:224] ^ 0);
  assign w908[22] = |(datain[223:220] ^ 11);
  assign w908[23] = |(datain[219:216] ^ 14);
  assign w908[24] = |(datain[215:212] ^ 0);
  assign w908[25] = |(datain[211:208] ^ 0);
  assign w908[26] = |(datain[207:204] ^ 0);
  assign w908[27] = |(datain[203:200] ^ 0);
  assign w908[28] = |(datain[199:196] ^ 1);
  assign w908[29] = |(datain[195:192] ^ 6);
  assign w908[30] = |(datain[191:188] ^ 1);
  assign w908[31] = |(datain[187:184] ^ 15);
  assign w908[32] = |(datain[183:180] ^ 11);
  assign w908[33] = |(datain[179:176] ^ 4);
  assign w908[34] = |(datain[175:172] ^ 4);
  assign w908[35] = |(datain[171:168] ^ 7);
  assign w908[36] = |(datain[167:164] ^ 12);
  assign w908[37] = |(datain[163:160] ^ 13);
  assign w908[38] = |(datain[159:156] ^ 2);
  assign w908[39] = |(datain[155:152] ^ 1);
  assign w908[40] = |(datain[151:148] ^ 0);
  assign w908[41] = |(datain[147:144] ^ 14);
  assign comp[908] = ~(|w908);
  wire [42-1:0] w909;
  assign w909[0] = |(datain[311:308] ^ 5);
  assign w909[1] = |(datain[307:304] ^ 13);
  assign w909[2] = |(datain[303:300] ^ 8);
  assign w909[3] = |(datain[299:296] ^ 3);
  assign w909[4] = |(datain[295:292] ^ 14);
  assign w909[5] = |(datain[291:288] ^ 13);
  assign w909[6] = |(datain[287:284] ^ 0);
  assign w909[7] = |(datain[283:280] ^ 3);
  assign w909[8] = |(datain[279:276] ^ 11);
  assign w909[9] = |(datain[275:272] ^ 9);
  assign w909[10] = |(datain[271:268] ^ 6);
  assign w909[11] = |(datain[267:264] ^ 1);
  assign w909[12] = |(datain[263:260] ^ 0);
  assign w909[13] = |(datain[259:256] ^ 3);
  assign w909[14] = |(datain[255:252] ^ 8);
  assign w909[15] = |(datain[251:248] ^ 11);
  assign w909[16] = |(datain[247:244] ^ 15);
  assign w909[17] = |(datain[243:240] ^ 13);
  assign w909[18] = |(datain[239:236] ^ 2);
  assign w909[19] = |(datain[235:232] ^ 14);
  assign w909[20] = |(datain[231:228] ^ 15);
  assign w909[21] = |(datain[227:224] ^ 6);
  assign w909[22] = |(datain[223:220] ^ 5);
  assign w909[23] = |(datain[219:216] ^ 5);
  assign w909[24] = |(datain[215:212] ^ 1);
  assign w909[25] = |(datain[211:208] ^ 3);
  assign w909[26] = |(datain[207:204] ^ 4);
  assign w909[27] = |(datain[203:200] ^ 7);
  assign w909[28] = |(datain[199:196] ^ 14);
  assign w909[29] = |(datain[195:192] ^ 2);
  assign w909[30] = |(datain[191:188] ^ 15);
  assign w909[31] = |(datain[187:184] ^ 9);
  assign w909[32] = |(datain[183:180] ^ 10);
  assign w909[33] = |(datain[179:176] ^ 15);
  assign w909[34] = |(datain[175:172] ^ 10);
  assign w909[35] = |(datain[171:168] ^ 13);
  assign w909[36] = |(datain[167:164] ^ 10);
  assign w909[37] = |(datain[163:160] ^ 9);
  assign w909[38] = |(datain[159:156] ^ 14);
  assign w909[39] = |(datain[155:152] ^ 1);
  assign w909[40] = |(datain[151:148] ^ 15);
  assign w909[41] = |(datain[147:144] ^ 9);
  assign comp[909] = ~(|w909);
  wire [44-1:0] w910;
  assign w910[0] = |(datain[311:308] ^ 9);
  assign w910[1] = |(datain[307:304] ^ 5);
  assign w910[2] = |(datain[303:300] ^ 11);
  assign w910[3] = |(datain[299:296] ^ 15);
  assign w910[4] = |(datain[295:292] ^ 12);
  assign w910[5] = |(datain[291:288] ^ 15);
  assign w910[6] = |(datain[287:284] ^ 0);
  assign w910[7] = |(datain[283:280] ^ 3);
  assign w910[8] = |(datain[279:276] ^ 0);
  assign w910[9] = |(datain[275:272] ^ 3);
  assign w910[10] = |(datain[271:268] ^ 15);
  assign w910[11] = |(datain[267:264] ^ 13);
  assign w910[12] = |(datain[263:260] ^ 2);
  assign w910[13] = |(datain[259:256] ^ 14);
  assign w910[14] = |(datain[255:252] ^ 8);
  assign w910[15] = |(datain[251:248] ^ 1);
  assign w910[16] = |(datain[247:244] ^ 3);
  assign w910[17] = |(datain[243:240] ^ 13);
  assign w910[18] = |(datain[239:236] ^ 12);
  assign w910[19] = |(datain[235:232] ^ 3);
  assign w910[20] = |(datain[231:228] ^ 12);
  assign w910[21] = |(datain[227:224] ^ 3);
  assign w910[22] = |(datain[223:220] ^ 7);
  assign w910[23] = |(datain[219:216] ^ 4);
  assign w910[24] = |(datain[215:212] ^ 1);
  assign w910[25] = |(datain[211:208] ^ 6);
  assign w910[26] = |(datain[207:204] ^ 11);
  assign w910[27] = |(datain[203:200] ^ 9);
  assign w910[28] = |(datain[199:196] ^ 11);
  assign w910[29] = |(datain[195:192] ^ 14);
  assign w910[30] = |(datain[191:188] ^ 0);
  assign w910[31] = |(datain[187:184] ^ 3);
  assign w910[32] = |(datain[183:180] ^ 11);
  assign w910[33] = |(datain[179:176] ^ 15);
  assign w910[34] = |(datain[175:172] ^ 2);
  assign w910[35] = |(datain[171:168] ^ 10);
  assign w910[36] = |(datain[167:164] ^ 0);
  assign w910[37] = |(datain[163:160] ^ 0);
  assign w910[38] = |(datain[159:156] ^ 0);
  assign w910[39] = |(datain[155:152] ^ 3);
  assign w910[40] = |(datain[151:148] ^ 15);
  assign w910[41] = |(datain[147:144] ^ 13);
  assign w910[42] = |(datain[143:140] ^ 11);
  assign w910[43] = |(datain[139:136] ^ 2);
  assign comp[910] = ~(|w910);
  wire [44-1:0] w911;
  assign w911[0] = |(datain[311:308] ^ 11);
  assign w911[1] = |(datain[307:304] ^ 15);
  assign w911[2] = |(datain[303:300] ^ 3);
  assign w911[3] = |(datain[299:296] ^ 9);
  assign w911[4] = |(datain[295:292] ^ 0);
  assign w911[5] = |(datain[291:288] ^ 0);
  assign w911[6] = |(datain[287:284] ^ 0);
  assign w911[7] = |(datain[283:280] ^ 3);
  assign w911[8] = |(datain[279:276] ^ 15);
  assign w911[9] = |(datain[275:272] ^ 13);
  assign w911[10] = |(datain[271:268] ^ 11);
  assign w911[11] = |(datain[267:264] ^ 2);
  assign w911[12] = |(datain[263:260] ^ 0);
  assign w911[13] = |(datain[259:256] ^ 1);
  assign w911[14] = |(datain[255:252] ^ 2);
  assign w911[15] = |(datain[251:248] ^ 14);
  assign w911[16] = |(datain[247:244] ^ 3);
  assign w911[17] = |(datain[243:240] ^ 0);
  assign w911[18] = |(datain[239:236] ^ 1);
  assign w911[19] = |(datain[235:232] ^ 5);
  assign w911[20] = |(datain[231:228] ^ 2);
  assign w911[21] = |(datain[227:224] ^ 14);
  assign w911[22] = |(datain[223:220] ^ 2);
  assign w911[23] = |(datain[219:216] ^ 8);
  assign w911[24] = |(datain[215:212] ^ 0);
  assign w911[25] = |(datain[211:208] ^ 13);
  assign w911[26] = |(datain[207:204] ^ 9);
  assign w911[27] = |(datain[203:200] ^ 0);
  assign w911[28] = |(datain[199:196] ^ 9);
  assign w911[29] = |(datain[195:192] ^ 0);
  assign w911[30] = |(datain[191:188] ^ 9);
  assign w911[31] = |(datain[187:184] ^ 0);
  assign w911[32] = |(datain[183:180] ^ 2);
  assign w911[33] = |(datain[179:176] ^ 14);
  assign w911[34] = |(datain[175:172] ^ 2);
  assign w911[35] = |(datain[171:168] ^ 8);
  assign w911[36] = |(datain[167:164] ^ 1);
  assign w911[37] = |(datain[163:160] ^ 5);
  assign w911[38] = |(datain[159:156] ^ 4);
  assign w911[39] = |(datain[155:152] ^ 7);
  assign w911[40] = |(datain[151:148] ^ 14);
  assign w911[41] = |(datain[147:144] ^ 2);
  assign w911[42] = |(datain[143:140] ^ 15);
  assign w911[43] = |(datain[139:136] ^ 1);
  assign comp[911] = ~(|w911);
  wire [74-1:0] w912;
  assign w912[0] = |(datain[311:308] ^ 7);
  assign w912[1] = |(datain[307:304] ^ 13);
  assign w912[2] = |(datain[303:300] ^ 0);
  assign w912[3] = |(datain[299:296] ^ 2);
  assign w912[4] = |(datain[295:292] ^ 4);
  assign w912[5] = |(datain[291:288] ^ 13);
  assign w912[6] = |(datain[287:284] ^ 7);
  assign w912[7] = |(datain[283:280] ^ 5);
  assign w912[8] = |(datain[279:276] ^ 0);
  assign w912[9] = |(datain[275:272] ^ 1);
  assign w912[10] = |(datain[271:268] ^ 15);
  assign w912[11] = |(datain[267:264] ^ 9);
  assign w912[12] = |(datain[263:260] ^ 12);
  assign w912[13] = |(datain[259:256] ^ 3);
  assign w912[14] = |(datain[255:252] ^ 5);
  assign w912[15] = |(datain[251:248] ^ 0);
  assign w912[16] = |(datain[247:244] ^ 5);
  assign w912[17] = |(datain[243:240] ^ 6);
  assign w912[18] = |(datain[239:236] ^ 5);
  assign w912[19] = |(datain[235:232] ^ 7);
  assign w912[20] = |(datain[231:228] ^ 5);
  assign w912[21] = |(datain[227:224] ^ 1);
  assign w912[22] = |(datain[223:220] ^ 5);
  assign w912[23] = |(datain[219:216] ^ 3);
  assign w912[24] = |(datain[215:212] ^ 1);
  assign w912[25] = |(datain[211:208] ^ 14);
  assign w912[26] = |(datain[207:204] ^ 0);
  assign w912[27] = |(datain[203:200] ^ 6);
  assign w912[28] = |(datain[199:196] ^ 9);
  assign w912[29] = |(datain[195:192] ^ 12);
  assign w912[30] = |(datain[191:188] ^ 11);
  assign w912[31] = |(datain[187:184] ^ 4);
  assign w912[32] = |(datain[183:180] ^ 6);
  assign w912[33] = |(datain[179:176] ^ 2);
  assign w912[34] = |(datain[175:172] ^ 12);
  assign w912[35] = |(datain[171:168] ^ 13);
  assign w912[36] = |(datain[167:164] ^ 2);
  assign w912[37] = |(datain[163:160] ^ 1);
  assign w912[38] = |(datain[159:156] ^ 5);
  assign w912[39] = |(datain[155:152] ^ 3);
  assign w912[40] = |(datain[151:148] ^ 1);
  assign w912[41] = |(datain[147:144] ^ 15);
  assign w912[42] = |(datain[143:140] ^ 10);
  assign w912[43] = |(datain[139:136] ^ 1);
  assign w912[44] = |(datain[135:132] ^ 2);
  assign w912[45] = |(datain[131:128] ^ 12);
  assign w912[46] = |(datain[127:124] ^ 0);
  assign w912[47] = |(datain[123:120] ^ 0);
  assign w912[48] = |(datain[119:116] ^ 5);
  assign w912[49] = |(datain[115:112] ^ 0);
  assign w912[50] = |(datain[111:108] ^ 1);
  assign w912[51] = |(datain[107:104] ^ 15);
  assign w912[52] = |(datain[103:100] ^ 3);
  assign w912[53] = |(datain[99:96] ^ 3);
  assign w912[54] = |(datain[95:92] ^ 15);
  assign w912[55] = |(datain[91:88] ^ 6);
  assign w912[56] = |(datain[87:84] ^ 4);
  assign w912[57] = |(datain[83:80] ^ 6);
  assign w912[58] = |(datain[79:76] ^ 8);
  assign w912[59] = |(datain[75:72] ^ 0);
  assign w912[60] = |(datain[71:68] ^ 3);
  assign w912[61] = |(datain[67:64] ^ 12);
  assign w912[62] = |(datain[63:60] ^ 0);
  assign w912[63] = |(datain[59:56] ^ 1);
  assign w912[64] = |(datain[55:52] ^ 7);
  assign w912[65] = |(datain[51:48] ^ 5);
  assign w912[66] = |(datain[47:44] ^ 15);
  assign w912[67] = |(datain[43:40] ^ 10);
  assign w912[68] = |(datain[39:36] ^ 4);
  assign w912[69] = |(datain[35:32] ^ 6);
  assign w912[70] = |(datain[31:28] ^ 4);
  assign w912[71] = |(datain[27:24] ^ 6);
  assign w912[72] = |(datain[23:20] ^ 4);
  assign w912[73] = |(datain[19:16] ^ 6);
  assign comp[912] = ~(|w912);
  wire [76-1:0] w913;
  assign w913[0] = |(datain[311:308] ^ 0);
  assign w913[1] = |(datain[307:304] ^ 7);
  assign w913[2] = |(datain[303:300] ^ 9);
  assign w913[3] = |(datain[299:296] ^ 0);
  assign w913[4] = |(datain[295:292] ^ 14);
  assign w913[5] = |(datain[291:288] ^ 8);
  assign w913[6] = |(datain[287:284] ^ 1);
  assign w913[7] = |(datain[283:280] ^ 7);
  assign w913[8] = |(datain[279:276] ^ 0);
  assign w913[9] = |(datain[275:272] ^ 2);
  assign w913[10] = |(datain[271:268] ^ 14);
  assign w913[11] = |(datain[267:264] ^ 11);
  assign w913[12] = |(datain[263:260] ^ 0);
  assign w913[13] = |(datain[259:256] ^ 8);
  assign w913[14] = |(datain[255:252] ^ 9);
  assign w913[15] = |(datain[251:248] ^ 0);
  assign w913[16] = |(datain[247:244] ^ 5);
  assign w913[17] = |(datain[243:240] ^ 11);
  assign w913[18] = |(datain[239:236] ^ 5);
  assign w913[19] = |(datain[235:232] ^ 9);
  assign w913[20] = |(datain[231:228] ^ 9);
  assign w913[21] = |(datain[227:224] ^ 13);
  assign w913[22] = |(datain[223:220] ^ 15);
  assign w913[23] = |(datain[219:216] ^ 9);
  assign w913[24] = |(datain[215:212] ^ 9);
  assign w913[25] = |(datain[211:208] ^ 12);
  assign w913[26] = |(datain[207:204] ^ 5);
  assign w913[27] = |(datain[203:200] ^ 1);
  assign w913[28] = |(datain[199:196] ^ 5);
  assign w913[29] = |(datain[195:192] ^ 3);
  assign w913[30] = |(datain[191:188] ^ 12);
  assign w913[31] = |(datain[187:184] ^ 15);
  assign w913[32] = |(datain[183:180] ^ 11);
  assign w913[33] = |(datain[179:176] ^ 0);
  assign w913[34] = |(datain[175:172] ^ 1);
  assign w913[35] = |(datain[171:168] ^ 3);
  assign w913[36] = |(datain[167:164] ^ 12);
  assign w913[37] = |(datain[163:160] ^ 13);
  assign w913[38] = |(datain[159:156] ^ 2);
  assign w913[39] = |(datain[155:152] ^ 1);
  assign w913[40] = |(datain[151:148] ^ 14);
  assign w913[41] = |(datain[147:144] ^ 8);
  assign w913[42] = |(datain[143:140] ^ 9);
  assign w913[43] = |(datain[139:136] ^ 6);
  assign w913[44] = |(datain[135:132] ^ 0);
  assign w913[45] = |(datain[131:128] ^ 1);
  assign w913[46] = |(datain[127:124] ^ 12);
  assign w913[47] = |(datain[123:120] ^ 15);
  assign w913[48] = |(datain[119:116] ^ 5);
  assign w913[49] = |(datain[115:112] ^ 1);
  assign w913[50] = |(datain[111:108] ^ 1);
  assign w913[51] = |(datain[107:104] ^ 14);
  assign w913[52] = |(datain[103:100] ^ 5);
  assign w913[53] = |(datain[99:96] ^ 2);
  assign w913[54] = |(datain[95:92] ^ 5);
  assign w913[55] = |(datain[91:88] ^ 0);
  assign w913[56] = |(datain[87:84] ^ 8);
  assign w913[57] = |(datain[83:80] ^ 3);
  assign w913[58] = |(datain[79:76] ^ 15);
  assign w913[59] = |(datain[75:72] ^ 11);
  assign w913[60] = |(datain[71:68] ^ 0);
  assign w913[61] = |(datain[67:64] ^ 1);
  assign w913[62] = |(datain[63:60] ^ 7);
  assign w913[63] = |(datain[59:56] ^ 4);
  assign w913[64] = |(datain[55:52] ^ 1);
  assign w913[65] = |(datain[51:48] ^ 13);
  assign w913[66] = |(datain[47:44] ^ 11);
  assign w913[67] = |(datain[43:40] ^ 4);
  assign w913[68] = |(datain[39:36] ^ 2);
  assign w913[69] = |(datain[35:32] ^ 12);
  assign w913[70] = |(datain[31:28] ^ 12);
  assign w913[71] = |(datain[27:24] ^ 13);
  assign w913[72] = |(datain[23:20] ^ 2);
  assign w913[73] = |(datain[19:16] ^ 1);
  assign w913[74] = |(datain[15:12] ^ 8);
  assign w913[75] = |(datain[11:8] ^ 0);
  assign comp[913] = ~(|w913);
  wire [30-1:0] w914;
  assign w914[0] = |(datain[311:308] ^ 11);
  assign w914[1] = |(datain[307:304] ^ 9);
  assign w914[2] = |(datain[303:300] ^ 2);
  assign w914[3] = |(datain[299:296] ^ 4);
  assign w914[4] = |(datain[295:292] ^ 0);
  assign w914[5] = |(datain[291:288] ^ 1);
  assign w914[6] = |(datain[287:284] ^ 3);
  assign w914[7] = |(datain[283:280] ^ 0);
  assign w914[8] = |(datain[279:276] ^ 2);
  assign w914[9] = |(datain[275:272] ^ 4);
  assign w914[10] = |(datain[271:268] ^ 4);
  assign w914[11] = |(datain[267:264] ^ 6);
  assign w914[12] = |(datain[263:260] ^ 14);
  assign w914[13] = |(datain[259:256] ^ 2);
  assign w914[14] = |(datain[255:252] ^ 15);
  assign w914[15] = |(datain[251:248] ^ 11);
  assign w914[16] = |(datain[247:244] ^ 5);
  assign w914[17] = |(datain[243:240] ^ 14);
  assign w914[18] = |(datain[239:236] ^ 12);
  assign w914[19] = |(datain[235:232] ^ 3);
  assign w914[20] = |(datain[231:228] ^ 14);
  assign w914[21] = |(datain[227:224] ^ 8);
  assign w914[22] = |(datain[223:220] ^ 0);
  assign w914[23] = |(datain[219:216] ^ 1);
  assign w914[24] = |(datain[215:212] ^ 0);
  assign w914[25] = |(datain[211:208] ^ 0);
  assign w914[26] = |(datain[207:204] ^ 12);
  assign w914[27] = |(datain[203:200] ^ 15);
  assign w914[28] = |(datain[199:196] ^ 5);
  assign w914[29] = |(datain[195:192] ^ 13);
  assign comp[914] = ~(|w914);
  wire [42-1:0] w915;
  assign w915[0] = |(datain[311:308] ^ 2);
  assign w915[1] = |(datain[307:304] ^ 0);
  assign w915[2] = |(datain[303:300] ^ 11);
  assign w915[3] = |(datain[299:296] ^ 8);
  assign w915[4] = |(datain[295:292] ^ 14);
  assign w915[5] = |(datain[291:288] ^ 0);
  assign w915[6] = |(datain[287:284] ^ 14);
  assign w915[7] = |(datain[283:280] ^ 0);
  assign w915[8] = |(datain[279:276] ^ 12);
  assign w915[9] = |(datain[275:272] ^ 13);
  assign w915[10] = |(datain[271:268] ^ 2);
  assign w915[11] = |(datain[267:264] ^ 1);
  assign w915[12] = |(datain[263:260] ^ 0);
  assign w915[13] = |(datain[259:256] ^ 12);
  assign w915[14] = |(datain[255:252] ^ 0);
  assign w915[15] = |(datain[251:248] ^ 0);
  assign w915[16] = |(datain[247:244] ^ 7);
  assign w915[17] = |(datain[243:240] ^ 4);
  assign w915[18] = |(datain[239:236] ^ 0);
  assign w915[19] = |(datain[235:232] ^ 2);
  assign w915[20] = |(datain[231:228] ^ 12);
  assign w915[21] = |(datain[227:224] ^ 13);
  assign w915[22] = |(datain[223:220] ^ 2);
  assign w915[23] = |(datain[219:216] ^ 0);
  assign w915[24] = |(datain[215:212] ^ 14);
  assign w915[25] = |(datain[211:208] ^ 4);
  assign w915[26] = |(datain[207:204] ^ 4);
  assign w915[27] = |(datain[203:200] ^ 0);
  assign w915[28] = |(datain[199:196] ^ 0);
  assign w915[29] = |(datain[195:192] ^ 10);
  assign w915[30] = |(datain[191:188] ^ 12);
  assign w915[31] = |(datain[187:184] ^ 0);
  assign w915[32] = |(datain[183:180] ^ 7);
  assign w915[33] = |(datain[179:176] ^ 5);
  assign w915[34] = |(datain[175:172] ^ 0);
  assign w915[35] = |(datain[171:168] ^ 2);
  assign w915[36] = |(datain[167:164] ^ 12);
  assign w915[37] = |(datain[163:160] ^ 13);
  assign w915[38] = |(datain[159:156] ^ 2);
  assign w915[39] = |(datain[155:152] ^ 0);
  assign w915[40] = |(datain[151:148] ^ 5);
  assign w915[41] = |(datain[147:144] ^ 8);
  assign comp[915] = ~(|w915);
  wire [30-1:0] w916;
  assign w916[0] = |(datain[311:308] ^ 13);
  assign w916[1] = |(datain[307:304] ^ 2);
  assign w916[2] = |(datain[303:300] ^ 11);
  assign w916[3] = |(datain[299:296] ^ 9);
  assign w916[4] = |(datain[295:292] ^ 0);
  assign w916[5] = |(datain[291:288] ^ 0);
  assign w916[6] = |(datain[287:284] ^ 14);
  assign w916[7] = |(datain[283:280] ^ 15);
  assign w916[8] = |(datain[279:276] ^ 11);
  assign w916[9] = |(datain[275:272] ^ 4);
  assign w916[10] = |(datain[271:268] ^ 3);
  assign w916[11] = |(datain[267:264] ^ 15);
  assign w916[12] = |(datain[263:260] ^ 9);
  assign w916[13] = |(datain[259:256] ^ 12);
  assign w916[14] = |(datain[255:252] ^ 15);
  assign w916[15] = |(datain[251:248] ^ 10);
  assign w916[16] = |(datain[247:244] ^ 0);
  assign w916[17] = |(datain[243:240] ^ 14);
  assign w916[18] = |(datain[239:236] ^ 14);
  assign w916[19] = |(datain[235:232] ^ 8);
  assign w916[20] = |(datain[231:228] ^ 0);
  assign w916[21] = |(datain[227:224] ^ 11);
  assign w916[22] = |(datain[223:220] ^ 0);
  assign w916[23] = |(datain[219:216] ^ 0);
  assign w916[24] = |(datain[215:212] ^ 12);
  assign w916[25] = |(datain[211:208] ^ 3);
  assign w916[26] = |(datain[207:204] ^ 3);
  assign w916[27] = |(datain[203:200] ^ 13);
  assign w916[28] = |(datain[199:196] ^ 0);
  assign w916[29] = |(datain[195:192] ^ 0);
  assign comp[916] = ~(|w916);
  wire [74-1:0] w917;
  assign w917[0] = |(datain[311:308] ^ 5);
  assign w917[1] = |(datain[307:304] ^ 0);
  assign w917[2] = |(datain[303:300] ^ 15);
  assign w917[3] = |(datain[299:296] ^ 12);
  assign w917[4] = |(datain[295:292] ^ 15);
  assign w917[5] = |(datain[291:288] ^ 3);
  assign w917[6] = |(datain[287:284] ^ 10);
  assign w917[7] = |(datain[283:280] ^ 4);
  assign w917[8] = |(datain[279:276] ^ 12);
  assign w917[9] = |(datain[275:272] ^ 11);
  assign w917[10] = |(datain[271:268] ^ 9);
  assign w917[11] = |(datain[267:264] ^ 9);
  assign w917[12] = |(datain[263:260] ^ 2);
  assign w917[13] = |(datain[259:256] ^ 11);
  assign w917[14] = |(datain[255:252] ^ 13);
  assign w917[15] = |(datain[251:248] ^ 11);
  assign w917[16] = |(datain[247:244] ^ 12);
  assign w917[17] = |(datain[243:240] ^ 13);
  assign w917[18] = |(datain[239:236] ^ 1);
  assign w917[19] = |(datain[235:232] ^ 3);
  assign w917[20] = |(datain[231:228] ^ 11);
  assign w917[21] = |(datain[227:224] ^ 8);
  assign w917[22] = |(datain[223:220] ^ 0);
  assign w917[23] = |(datain[219:216] ^ 15);
  assign w917[24] = |(datain[215:212] ^ 0);
  assign w917[25] = |(datain[211:208] ^ 5);
  assign w917[26] = |(datain[207:204] ^ 8);
  assign w917[27] = |(datain[203:200] ^ 4);
  assign w917[28] = |(datain[199:196] ^ 0);
  assign w917[29] = |(datain[195:192] ^ 6);
  assign w917[30] = |(datain[191:188] ^ 6);
  assign w917[31] = |(datain[187:184] ^ 12);
  assign w917[32] = |(datain[183:180] ^ 0);
  assign w917[33] = |(datain[179:176] ^ 4);
  assign w917[34] = |(datain[175:172] ^ 7);
  assign w917[35] = |(datain[171:168] ^ 5);
  assign w917[36] = |(datain[167:164] ^ 0);
  assign w917[37] = |(datain[163:160] ^ 3);
  assign w917[38] = |(datain[159:156] ^ 4);
  assign w917[39] = |(datain[155:152] ^ 1);
  assign w917[40] = |(datain[151:148] ^ 12);
  assign w917[41] = |(datain[147:144] ^ 13);
  assign w917[42] = |(datain[143:140] ^ 1);
  assign w917[43] = |(datain[139:136] ^ 3);
  assign w917[44] = |(datain[135:132] ^ 11);
  assign w917[45] = |(datain[131:128] ^ 2);
  assign w917[46] = |(datain[127:124] ^ 8);
  assign w917[47] = |(datain[123:120] ^ 0);
  assign w917[48] = |(datain[119:116] ^ 5);
  assign w917[49] = |(datain[115:112] ^ 2);
  assign w917[50] = |(datain[111:108] ^ 0);
  assign w917[51] = |(datain[107:104] ^ 14);
  assign w917[52] = |(datain[103:100] ^ 1);
  assign w917[53] = |(datain[99:96] ^ 15);
  assign w917[54] = |(datain[95:92] ^ 11);
  assign w917[55] = |(datain[91:88] ^ 4);
  assign w917[56] = |(datain[87:84] ^ 0);
  assign w917[57] = |(datain[83:80] ^ 8);
  assign w917[58] = |(datain[79:76] ^ 12);
  assign w917[59] = |(datain[75:72] ^ 13);
  assign w917[60] = |(datain[71:68] ^ 1);
  assign w917[61] = |(datain[67:64] ^ 3);
  assign w917[62] = |(datain[63:60] ^ 8);
  assign w917[63] = |(datain[59:56] ^ 8);
  assign w917[64] = |(datain[55:52] ^ 7);
  assign w917[65] = |(datain[51:48] ^ 5);
  assign w917[66] = |(datain[47:44] ^ 12);
  assign w917[67] = |(datain[43:40] ^ 8);
  assign w917[68] = |(datain[39:36] ^ 8);
  assign w917[69] = |(datain[35:32] ^ 3);
  assign w917[70] = |(datain[31:28] ^ 14);
  assign w917[71] = |(datain[27:24] ^ 1);
  assign w917[72] = |(datain[23:20] ^ 3);
  assign w917[73] = |(datain[19:16] ^ 15);
  assign comp[917] = ~(|w917);
  wire [38-1:0] w918;
  assign w918[0] = |(datain[311:308] ^ 8);
  assign w918[1] = |(datain[307:304] ^ 14);
  assign w918[2] = |(datain[303:300] ^ 12);
  assign w918[3] = |(datain[299:296] ^ 0);
  assign w918[4] = |(datain[295:292] ^ 11);
  assign w918[5] = |(datain[291:288] ^ 8);
  assign w918[6] = |(datain[287:284] ^ 0);
  assign w918[7] = |(datain[283:280] ^ 1);
  assign w918[8] = |(datain[279:276] ^ 0);
  assign w918[9] = |(datain[275:272] ^ 2);
  assign w918[10] = |(datain[271:268] ^ 11);
  assign w918[11] = |(datain[267:264] ^ 11);
  assign w918[12] = |(datain[263:260] ^ 0);
  assign w918[13] = |(datain[259:256] ^ 0);
  assign w918[14] = |(datain[255:252] ^ 0);
  assign w918[15] = |(datain[251:248] ^ 8);
  assign w918[16] = |(datain[247:244] ^ 11);
  assign w918[17] = |(datain[243:240] ^ 9);
  assign w918[18] = |(datain[239:236] ^ 0);
  assign w918[19] = |(datain[235:232] ^ 0);
  assign w918[20] = |(datain[231:228] ^ 0);
  assign w918[21] = |(datain[227:224] ^ 0);
  assign w918[22] = |(datain[223:220] ^ 11);
  assign w918[23] = |(datain[219:216] ^ 6);
  assign w918[24] = |(datain[215:212] ^ 0);
  assign w918[25] = |(datain[211:208] ^ 0);
  assign w918[26] = |(datain[207:204] ^ 12);
  assign w918[27] = |(datain[203:200] ^ 13);
  assign w918[28] = |(datain[199:196] ^ 1);
  assign w918[29] = |(datain[195:192] ^ 3);
  assign w918[30] = |(datain[191:188] ^ 14);
  assign w918[31] = |(datain[187:184] ^ 10);
  assign w918[32] = |(datain[183:180] ^ 7);
  assign w918[33] = |(datain[179:176] ^ 0);
  assign w918[34] = |(datain[175:172] ^ 0);
  assign w918[35] = |(datain[171:168] ^ 8);
  assign w918[36] = |(datain[167:164] ^ 0);
  assign w918[37] = |(datain[163:160] ^ 0);
  assign comp[918] = ~(|w918);
  wire [74-1:0] w919;
  assign w919[0] = |(datain[311:308] ^ 5);
  assign w919[1] = |(datain[307:304] ^ 0);
  assign w919[2] = |(datain[303:300] ^ 12);
  assign w919[3] = |(datain[299:296] ^ 11);
  assign w919[4] = |(datain[295:292] ^ 11);
  assign w919[5] = |(datain[291:288] ^ 15);
  assign w919[6] = |(datain[287:284] ^ 12);
  assign w919[7] = |(datain[283:280] ^ 0);
  assign w919[8] = |(datain[279:276] ^ 0);
  assign w919[9] = |(datain[275:272] ^ 0);
  assign w919[10] = |(datain[271:268] ^ 14);
  assign w919[11] = |(datain[267:264] ^ 8);
  assign w919[12] = |(datain[263:260] ^ 4);
  assign w919[13] = |(datain[259:256] ^ 5);
  assign w919[14] = |(datain[255:252] ^ 0);
  assign w919[15] = |(datain[251:248] ^ 0);
  assign w919[16] = |(datain[247:244] ^ 3);
  assign w919[17] = |(datain[243:240] ^ 3);
  assign w919[18] = |(datain[239:236] ^ 12);
  assign w919[19] = |(datain[235:232] ^ 0);
  assign w919[20] = |(datain[231:228] ^ 12);
  assign w919[21] = |(datain[227:224] ^ 13);
  assign w919[22] = |(datain[223:220] ^ 1);
  assign w919[23] = |(datain[219:216] ^ 10);
  assign w919[24] = |(datain[215:212] ^ 8);
  assign w919[25] = |(datain[211:208] ^ 1);
  assign w919[26] = |(datain[207:204] ^ 12);
  assign w919[27] = |(datain[203:200] ^ 2);
  assign w919[28] = |(datain[199:196] ^ 2);
  assign w919[29] = |(datain[195:192] ^ 2);
  assign w919[30] = |(datain[191:188] ^ 0);
  assign w919[31] = |(datain[187:184] ^ 2);
  assign w919[32] = |(datain[183:180] ^ 8);
  assign w919[33] = |(datain[179:176] ^ 3);
  assign w919[34] = |(datain[175:172] ^ 13);
  assign w919[35] = |(datain[171:168] ^ 1);
  assign w919[36] = |(datain[167:164] ^ 0);
  assign w919[37] = |(datain[163:160] ^ 0);
  assign w919[38] = |(datain[159:156] ^ 8);
  assign w919[39] = |(datain[155:152] ^ 11);
  assign w919[40] = |(datain[151:148] ^ 15);
  assign w919[41] = |(datain[147:144] ^ 2);
  assign w919[42] = |(datain[143:140] ^ 8);
  assign w919[43] = |(datain[139:136] ^ 11);
  assign w919[44] = |(datain[135:132] ^ 15);
  assign w919[45] = |(datain[131:128] ^ 9);
  assign w919[46] = |(datain[127:124] ^ 3);
  assign w919[47] = |(datain[123:120] ^ 3);
  assign w919[48] = |(datain[119:116] ^ 12);
  assign w919[49] = |(datain[115:112] ^ 0);
  assign w919[50] = |(datain[111:108] ^ 12);
  assign w919[51] = |(datain[107:104] ^ 13);
  assign w919[52] = |(datain[103:100] ^ 1);
  assign w919[53] = |(datain[99:96] ^ 10);
  assign w919[54] = |(datain[95:92] ^ 3);
  assign w919[55] = |(datain[91:88] ^ 11);
  assign w919[56] = |(datain[87:84] ^ 12);
  assign w919[57] = |(datain[83:80] ^ 15);
  assign w919[58] = |(datain[79:76] ^ 7);
  assign w919[59] = |(datain[75:72] ^ 12);
  assign w919[60] = |(datain[71:68] ^ 15);
  assign w919[61] = |(datain[67:64] ^ 8);
  assign w919[62] = |(datain[63:60] ^ 7);
  assign w919[63] = |(datain[59:56] ^ 7);
  assign w919[64] = |(datain[55:52] ^ 0);
  assign w919[65] = |(datain[51:48] ^ 4);
  assign w919[66] = |(datain[47:44] ^ 3);
  assign w919[67] = |(datain[43:40] ^ 11);
  assign w919[68] = |(datain[39:36] ^ 13);
  assign w919[69] = |(datain[35:32] ^ 6);
  assign w919[70] = |(datain[31:28] ^ 7);
  assign w919[71] = |(datain[27:24] ^ 12);
  assign w919[72] = |(datain[23:20] ^ 15);
  assign w919[73] = |(datain[19:16] ^ 2);
  assign comp[919] = ~(|w919);
  wire [74-1:0] w920;
  assign w920[0] = |(datain[311:308] ^ 3);
  assign w920[1] = |(datain[307:304] ^ 3);
  assign w920[2] = |(datain[303:300] ^ 15);
  assign w920[3] = |(datain[299:296] ^ 15);
  assign w920[4] = |(datain[295:292] ^ 15);
  assign w920[5] = |(datain[291:288] ^ 10);
  assign w920[6] = |(datain[287:284] ^ 8);
  assign w920[7] = |(datain[283:280] ^ 14);
  assign w920[8] = |(datain[279:276] ^ 13);
  assign w920[9] = |(datain[275:272] ^ 7);
  assign w920[10] = |(datain[271:268] ^ 8);
  assign w920[11] = |(datain[267:264] ^ 11);
  assign w920[12] = |(datain[263:260] ^ 14);
  assign w920[13] = |(datain[259:256] ^ 6);
  assign w920[14] = |(datain[255:252] ^ 15);
  assign w920[15] = |(datain[251:248] ^ 11);
  assign w920[16] = |(datain[247:244] ^ 8);
  assign w920[17] = |(datain[243:240] ^ 14);
  assign w920[18] = |(datain[239:236] ^ 13);
  assign w920[19] = |(datain[235:232] ^ 15);
  assign w920[20] = |(datain[231:228] ^ 12);
  assign w920[21] = |(datain[227:224] ^ 13);
  assign w920[22] = |(datain[223:220] ^ 1);
  assign w920[23] = |(datain[219:216] ^ 2);
  assign w920[24] = |(datain[215:212] ^ 4);
  assign w920[25] = |(datain[211:208] ^ 8);
  assign w920[26] = |(datain[207:204] ^ 10);
  assign w920[27] = |(datain[203:200] ^ 3);
  assign w920[28] = |(datain[199:196] ^ 1);
  assign w920[29] = |(datain[195:192] ^ 3);
  assign w920[30] = |(datain[191:188] ^ 0);
  assign w920[31] = |(datain[187:184] ^ 4);
  assign w920[32] = |(datain[183:180] ^ 12);
  assign w920[33] = |(datain[179:176] ^ 1);
  assign w920[34] = |(datain[175:172] ^ 14);
  assign w920[35] = |(datain[171:168] ^ 0);
  assign w920[36] = |(datain[167:164] ^ 0);
  assign w920[37] = |(datain[163:160] ^ 6);
  assign w920[38] = |(datain[159:156] ^ 8);
  assign w920[39] = |(datain[155:152] ^ 14);
  assign w920[40] = |(datain[151:148] ^ 12);
  assign w920[41] = |(datain[147:144] ^ 0);
  assign w920[42] = |(datain[143:140] ^ 15);
  assign w920[43] = |(datain[139:136] ^ 12);
  assign w920[44] = |(datain[135:132] ^ 11);
  assign w920[45] = |(datain[131:128] ^ 9);
  assign w920[46] = |(datain[127:124] ^ 0);
  assign w920[47] = |(datain[123:120] ^ 0);
  assign w920[48] = |(datain[119:116] ^ 0);
  assign w920[49] = |(datain[115:112] ^ 1);
  assign w920[50] = |(datain[111:108] ^ 15);
  assign w920[51] = |(datain[107:104] ^ 3);
  assign w920[52] = |(datain[103:100] ^ 10);
  assign w920[53] = |(datain[99:96] ^ 5);
  assign w920[54] = |(datain[95:92] ^ 0);
  assign w920[55] = |(datain[91:88] ^ 6);
  assign w920[56] = |(datain[87:84] ^ 6);
  assign w920[57] = |(datain[83:80] ^ 8);
  assign w920[58] = |(datain[79:76] ^ 6);
  assign w920[59] = |(datain[75:72] ^ 1);
  assign w920[60] = |(datain[71:68] ^ 0);
  assign w920[61] = |(datain[67:64] ^ 0);
  assign w920[62] = |(datain[63:60] ^ 12);
  assign w920[63] = |(datain[59:56] ^ 11);
  assign w920[64] = |(datain[55:52] ^ 14);
  assign w920[65] = |(datain[51:48] ^ 8);
  assign w920[66] = |(datain[47:44] ^ 5);
  assign w920[67] = |(datain[43:40] ^ 0);
  assign w920[68] = |(datain[39:36] ^ 0);
  assign w920[69] = |(datain[35:32] ^ 1);
  assign w920[70] = |(datain[31:28] ^ 12);
  assign w920[71] = |(datain[27:24] ^ 13);
  assign w920[72] = |(datain[23:20] ^ 1);
  assign w920[73] = |(datain[19:16] ^ 9);
  assign comp[920] = ~(|w920);
  wire [74-1:0] w921;
  assign w921[0] = |(datain[311:308] ^ 11);
  assign w921[1] = |(datain[307:304] ^ 8);
  assign w921[2] = |(datain[303:300] ^ 0);
  assign w921[3] = |(datain[299:296] ^ 1);
  assign w921[4] = |(datain[295:292] ^ 0);
  assign w921[5] = |(datain[291:288] ^ 3);
  assign w921[6] = |(datain[287:284] ^ 3);
  assign w921[7] = |(datain[283:280] ^ 3);
  assign w921[8] = |(datain[279:276] ^ 13);
  assign w921[9] = |(datain[275:272] ^ 11);
  assign w921[10] = |(datain[271:268] ^ 12);
  assign w921[11] = |(datain[267:264] ^ 13);
  assign w921[12] = |(datain[263:260] ^ 1);
  assign w921[13] = |(datain[259:256] ^ 3);
  assign w921[14] = |(datain[255:252] ^ 3);
  assign w921[15] = |(datain[251:248] ^ 2);
  assign w921[16] = |(datain[247:244] ^ 15);
  assign w921[17] = |(datain[243:240] ^ 6);
  assign w921[18] = |(datain[239:236] ^ 11);
  assign w921[19] = |(datain[235:232] ^ 9);
  assign w921[20] = |(datain[231:228] ^ 0);
  assign w921[21] = |(datain[227:224] ^ 13);
  assign w921[22] = |(datain[223:220] ^ 0);
  assign w921[23] = |(datain[219:216] ^ 0);
  assign w921[24] = |(datain[215:212] ^ 11);
  assign w921[25] = |(datain[211:208] ^ 11);
  assign w921[26] = |(datain[207:204] ^ 0);
  assign w921[27] = |(datain[203:200] ^ 0);
  assign w921[28] = |(datain[199:196] ^ 0);
  assign w921[29] = |(datain[195:192] ^ 2);
  assign w921[30] = |(datain[191:188] ^ 11);
  assign w921[31] = |(datain[187:184] ^ 8);
  assign w921[32] = |(datain[183:180] ^ 0);
  assign w921[33] = |(datain[179:176] ^ 1);
  assign w921[34] = |(datain[175:172] ^ 0);
  assign w921[35] = |(datain[171:168] ^ 3);
  assign w921[36] = |(datain[167:164] ^ 12);
  assign w921[37] = |(datain[163:160] ^ 13);
  assign w921[38] = |(datain[159:156] ^ 1);
  assign w921[39] = |(datain[155:152] ^ 3);
  assign w921[40] = |(datain[151:148] ^ 14);
  assign w921[41] = |(datain[147:144] ^ 8);
  assign w921[42] = |(datain[143:140] ^ 10);
  assign w921[43] = |(datain[139:136] ^ 7);
  assign w921[44] = |(datain[135:132] ^ 0);
  assign w921[45] = |(datain[131:128] ^ 0);
  assign w921[46] = |(datain[127:124] ^ 3);
  assign w921[47] = |(datain[123:120] ^ 2);
  assign w921[48] = |(datain[119:116] ^ 13);
  assign w921[49] = |(datain[115:112] ^ 2);
  assign w921[50] = |(datain[111:108] ^ 11);
  assign w921[51] = |(datain[107:104] ^ 8);
  assign w921[52] = |(datain[103:100] ^ 0);
  assign w921[53] = |(datain[99:96] ^ 1);
  assign w921[54] = |(datain[95:92] ^ 0);
  assign w921[55] = |(datain[91:88] ^ 2);
  assign w921[56] = |(datain[87:84] ^ 3);
  assign w921[57] = |(datain[83:80] ^ 3);
  assign w921[58] = |(datain[79:76] ^ 13);
  assign w921[59] = |(datain[75:72] ^ 11);
  assign w921[60] = |(datain[71:68] ^ 8);
  assign w921[61] = |(datain[67:64] ^ 14);
  assign w921[62] = |(datain[63:60] ^ 12);
  assign w921[63] = |(datain[59:56] ^ 3);
  assign w921[64] = |(datain[55:52] ^ 11);
  assign w921[65] = |(datain[51:48] ^ 11);
  assign w921[66] = |(datain[47:44] ^ 0);
  assign w921[67] = |(datain[43:40] ^ 0);
  assign w921[68] = |(datain[39:36] ^ 7);
  assign w921[69] = |(datain[35:32] ^ 12);
  assign w921[70] = |(datain[31:28] ^ 12);
  assign w921[71] = |(datain[27:24] ^ 13);
  assign w921[72] = |(datain[23:20] ^ 1);
  assign w921[73] = |(datain[19:16] ^ 3);
  assign comp[921] = ~(|w921);
  wire [76-1:0] w922;
  assign w922[0] = |(datain[311:308] ^ 8);
  assign w922[1] = |(datain[307:304] ^ 3);
  assign w922[2] = |(datain[303:300] ^ 12);
  assign w922[3] = |(datain[299:296] ^ 6);
  assign w922[4] = |(datain[295:292] ^ 0);
  assign w922[5] = |(datain[291:288] ^ 3);
  assign w922[6] = |(datain[287:284] ^ 11);
  assign w922[7] = |(datain[283:280] ^ 11);
  assign w922[8] = |(datain[279:276] ^ 0);
  assign w922[9] = |(datain[275:272] ^ 0);
  assign w922[10] = |(datain[271:268] ^ 7);
  assign w922[11] = |(datain[267:264] ^ 12);
  assign w922[12] = |(datain[263:260] ^ 8);
  assign w922[13] = |(datain[259:256] ^ 11);
  assign w922[14] = |(datain[255:252] ^ 15);
  assign w922[15] = |(datain[251:248] ^ 11);
  assign w922[16] = |(datain[247:244] ^ 8);
  assign w922[17] = |(datain[243:240] ^ 3);
  assign w922[18] = |(datain[239:236] ^ 12);
  assign w922[19] = |(datain[235:232] ^ 7);
  assign w922[20] = |(datain[231:228] ^ 0);
  assign w922[21] = |(datain[227:224] ^ 3);
  assign w922[22] = |(datain[223:220] ^ 0);
  assign w922[23] = |(datain[219:216] ^ 14);
  assign w922[24] = |(datain[215:212] ^ 0);
  assign w922[25] = |(datain[211:208] ^ 7);
  assign w922[26] = |(datain[207:204] ^ 15);
  assign w922[27] = |(datain[203:200] ^ 12);
  assign w922[28] = |(datain[199:196] ^ 15);
  assign w922[29] = |(datain[195:192] ^ 3);
  assign w922[30] = |(datain[191:188] ^ 10);
  assign w922[31] = |(datain[187:184] ^ 4);
  assign w922[32] = |(datain[183:180] ^ 8);
  assign w922[33] = |(datain[179:176] ^ 1);
  assign w922[34] = |(datain[175:172] ^ 12);
  assign w922[35] = |(datain[171:168] ^ 6);
  assign w922[36] = |(datain[167:164] ^ 9);
  assign w922[37] = |(datain[163:160] ^ 13);
  assign w922[38] = |(datain[159:156] ^ 0);
  assign w922[39] = |(datain[155:152] ^ 1);
  assign w922[40] = |(datain[151:148] ^ 8);
  assign w922[41] = |(datain[147:144] ^ 1);
  assign w922[42] = |(datain[143:140] ^ 12);
  assign w922[43] = |(datain[139:136] ^ 7);
  assign w922[44] = |(datain[135:132] ^ 9);
  assign w922[45] = |(datain[131:128] ^ 13);
  assign w922[46] = |(datain[127:124] ^ 0);
  assign w922[47] = |(datain[123:120] ^ 1);
  assign w922[48] = |(datain[119:116] ^ 11);
  assign w922[49] = |(datain[115:112] ^ 9);
  assign w922[50] = |(datain[111:108] ^ 3);
  assign w922[51] = |(datain[107:104] ^ 0);
  assign w922[52] = |(datain[103:100] ^ 0);
  assign w922[53] = |(datain[99:96] ^ 0);
  assign w922[54] = |(datain[95:92] ^ 15);
  assign w922[55] = |(datain[91:88] ^ 3);
  assign w922[56] = |(datain[87:84] ^ 10);
  assign w922[57] = |(datain[83:80] ^ 5);
  assign w922[58] = |(datain[79:76] ^ 8);
  assign w922[59] = |(datain[75:72] ^ 11);
  assign w922[60] = |(datain[71:68] ^ 13);
  assign w922[61] = |(datain[67:64] ^ 1);
  assign w922[62] = |(datain[63:60] ^ 4);
  assign w922[63] = |(datain[59:56] ^ 1);
  assign w922[64] = |(datain[55:52] ^ 11);
  assign w922[65] = |(datain[51:48] ^ 8);
  assign w922[66] = |(datain[47:44] ^ 0);
  assign w922[67] = |(datain[43:40] ^ 1);
  assign w922[68] = |(datain[39:36] ^ 0);
  assign w922[69] = |(datain[35:32] ^ 3);
  assign w922[70] = |(datain[31:28] ^ 12);
  assign w922[71] = |(datain[27:24] ^ 13);
  assign w922[72] = |(datain[23:20] ^ 13);
  assign w922[73] = |(datain[19:16] ^ 3);
  assign w922[74] = |(datain[15:12] ^ 5);
  assign w922[75] = |(datain[11:8] ^ 15);
  assign comp[922] = ~(|w922);
  wire [76-1:0] w923;
  assign w923[0] = |(datain[311:308] ^ 12);
  assign w923[1] = |(datain[307:304] ^ 13);
  assign w923[2] = |(datain[303:300] ^ 2);
  assign w923[3] = |(datain[299:296] ^ 15);
  assign w923[4] = |(datain[295:292] ^ 2);
  assign w923[5] = |(datain[291:288] ^ 14);
  assign w923[6] = |(datain[287:284] ^ 8);
  assign w923[7] = |(datain[283:280] ^ 12);
  assign w923[8] = |(datain[279:276] ^ 1);
  assign w923[9] = |(datain[275:272] ^ 14);
  assign w923[10] = |(datain[271:268] ^ 11);
  assign w923[11] = |(datain[267:264] ^ 8);
  assign w923[12] = |(datain[263:260] ^ 0);
  assign w923[13] = |(datain[259:256] ^ 1);
  assign w923[14] = |(datain[255:252] ^ 8);
  assign w923[15] = |(datain[251:248] ^ 11);
  assign w923[16] = |(datain[247:244] ^ 12);
  assign w923[17] = |(datain[243:240] ^ 10);
  assign w923[18] = |(datain[239:236] ^ 12);
  assign w923[19] = |(datain[235:232] ^ 13);
  assign w923[20] = |(datain[231:228] ^ 2);
  assign w923[21] = |(datain[227:224] ^ 15);
  assign w923[22] = |(datain[223:220] ^ 8);
  assign w923[23] = |(datain[219:216] ^ 9);
  assign w923[24] = |(datain[215:212] ^ 0);
  assign w923[25] = |(datain[211:208] ^ 14);
  assign w923[26] = |(datain[207:204] ^ 11);
  assign w923[27] = |(datain[203:200] ^ 6);
  assign w923[28] = |(datain[199:196] ^ 0);
  assign w923[29] = |(datain[195:192] ^ 1);
  assign w923[30] = |(datain[191:188] ^ 8);
  assign w923[31] = |(datain[187:184] ^ 0);
  assign w923[32] = |(datain[183:180] ^ 15);
  assign w923[33] = |(datain[179:176] ^ 9);
  assign w923[34] = |(datain[175:172] ^ 3);
  assign w923[35] = |(datain[171:168] ^ 2);
  assign w923[36] = |(datain[167:164] ^ 7);
  assign w923[37] = |(datain[163:160] ^ 4);
  assign w923[38] = |(datain[159:156] ^ 0);
  assign w923[39] = |(datain[155:152] ^ 10);
  assign w923[40] = |(datain[151:148] ^ 8);
  assign w923[41] = |(datain[147:144] ^ 12);
  assign w923[42] = |(datain[143:140] ^ 12);
  assign w923[43] = |(datain[139:136] ^ 9);
  assign w923[44] = |(datain[135:132] ^ 8);
  assign w923[45] = |(datain[131:128] ^ 3);
  assign w923[46] = |(datain[127:124] ^ 12);
  assign w923[47] = |(datain[123:120] ^ 1);
  assign w923[48] = |(datain[119:116] ^ 1);
  assign w923[49] = |(datain[115:112] ^ 0);
  assign w923[50] = |(datain[111:108] ^ 5);
  assign w923[51] = |(datain[107:104] ^ 1);
  assign w923[52] = |(datain[103:100] ^ 11);
  assign w923[53] = |(datain[99:96] ^ 8);
  assign w923[54] = |(datain[95:92] ^ 15);
  assign w923[55] = |(datain[91:88] ^ 13);
  assign w923[56] = |(datain[87:84] ^ 0);
  assign w923[57] = |(datain[83:80] ^ 0);
  assign w923[58] = |(datain[79:76] ^ 5);
  assign w923[59] = |(datain[75:72] ^ 0);
  assign w923[60] = |(datain[71:68] ^ 12);
  assign w923[61] = |(datain[67:64] ^ 11);
  assign w923[62] = |(datain[63:60] ^ 14);
  assign w923[63] = |(datain[59:56] ^ 8);
  assign w923[64] = |(datain[55:52] ^ 6);
  assign w923[65] = |(datain[51:48] ^ 8);
  assign w923[66] = |(datain[47:44] ^ 0);
  assign w923[67] = |(datain[43:40] ^ 0);
  assign w923[68] = |(datain[39:36] ^ 11);
  assign w923[69] = |(datain[35:32] ^ 4);
  assign w923[70] = |(datain[31:28] ^ 0);
  assign w923[71] = |(datain[27:24] ^ 4);
  assign w923[72] = |(datain[23:20] ^ 12);
  assign w923[73] = |(datain[19:16] ^ 13);
  assign w923[74] = |(datain[15:12] ^ 1);
  assign w923[75] = |(datain[11:8] ^ 10);
  assign comp[923] = ~(|w923);
  wire [76-1:0] w924;
  assign w924[0] = |(datain[311:308] ^ 0);
  assign w924[1] = |(datain[307:304] ^ 2);
  assign w924[2] = |(datain[303:300] ^ 11);
  assign w924[3] = |(datain[299:296] ^ 11);
  assign w924[4] = |(datain[295:292] ^ 0);
  assign w924[5] = |(datain[291:288] ^ 0);
  assign w924[6] = |(datain[287:284] ^ 0);
  assign w924[7] = |(datain[283:280] ^ 1);
  assign w924[8] = |(datain[279:276] ^ 5);
  assign w924[9] = |(datain[275:272] ^ 3);
  assign w924[10] = |(datain[271:268] ^ 2);
  assign w924[11] = |(datain[267:264] ^ 6);
  assign w924[12] = |(datain[263:260] ^ 8);
  assign w924[13] = |(datain[259:256] ^ 1);
  assign w924[14] = |(datain[255:252] ^ 3);
  assign w924[15] = |(datain[251:248] ^ 15);
  assign w924[16] = |(datain[247:244] ^ 5);
  assign w924[17] = |(datain[243:240] ^ 2);
  assign w924[18] = |(datain[239:236] ^ 2);
  assign w924[19] = |(datain[235:232] ^ 4);
  assign w924[20] = |(datain[231:228] ^ 7);
  assign w924[21] = |(datain[227:224] ^ 4);
  assign w924[22] = |(datain[223:220] ^ 0);
  assign w924[23] = |(datain[219:216] ^ 11);
  assign w924[24] = |(datain[215:212] ^ 12);
  assign w924[25] = |(datain[211:208] ^ 13);
  assign w924[26] = |(datain[207:204] ^ 1);
  assign w924[27] = |(datain[203:200] ^ 3);
  assign w924[28] = |(datain[199:196] ^ 5);
  assign w924[29] = |(datain[195:192] ^ 11);
  assign w924[30] = |(datain[191:188] ^ 7);
  assign w924[31] = |(datain[187:184] ^ 2);
  assign w924[32] = |(datain[183:180] ^ 1);
  assign w924[33] = |(datain[179:176] ^ 8);
  assign w924[34] = |(datain[175:172] ^ 0);
  assign w924[35] = |(datain[171:168] ^ 6);
  assign w924[36] = |(datain[167:164] ^ 11);
  assign w924[37] = |(datain[163:160] ^ 8);
  assign w924[38] = |(datain[159:156] ^ 0);
  assign w924[39] = |(datain[155:152] ^ 2);
  assign w924[40] = |(datain[151:148] ^ 0);
  assign w924[41] = |(datain[147:144] ^ 1);
  assign w924[42] = |(datain[143:140] ^ 5);
  assign w924[43] = |(datain[139:136] ^ 0);
  assign w924[44] = |(datain[135:132] ^ 12);
  assign w924[45] = |(datain[131:128] ^ 11);
  assign w924[46] = |(datain[127:124] ^ 11);
  assign w924[47] = |(datain[123:120] ^ 11);
  assign w924[48] = |(datain[119:116] ^ 0);
  assign w924[49] = |(datain[115:112] ^ 0);
  assign w924[50] = |(datain[111:108] ^ 0);
  assign w924[51] = |(datain[107:104] ^ 15);
  assign w924[52] = |(datain[103:100] ^ 11);
  assign w924[53] = |(datain[99:96] ^ 0);
  assign w924[54] = |(datain[95:92] ^ 0);
  assign w924[55] = |(datain[91:88] ^ 1);
  assign w924[56] = |(datain[87:84] ^ 11);
  assign w924[57] = |(datain[83:80] ^ 1);
  assign w924[58] = |(datain[79:76] ^ 0);
  assign w924[59] = |(datain[75:72] ^ 9);
  assign w924[60] = |(datain[71:68] ^ 12);
  assign w924[61] = |(datain[67:64] ^ 13);
  assign w924[62] = |(datain[63:60] ^ 1);
  assign w924[63] = |(datain[59:56] ^ 3);
  assign w924[64] = |(datain[55:52] ^ 5);
  assign w924[65] = |(datain[51:48] ^ 11);
  assign w924[66] = |(datain[47:44] ^ 7);
  assign w924[67] = |(datain[43:40] ^ 2);
  assign w924[68] = |(datain[39:36] ^ 0);
  assign w924[69] = |(datain[35:32] ^ 6);
  assign w924[70] = |(datain[31:28] ^ 0);
  assign w924[71] = |(datain[27:24] ^ 6);
  assign w924[72] = |(datain[23:20] ^ 11);
  assign w924[73] = |(datain[19:16] ^ 8);
  assign w924[74] = |(datain[15:12] ^ 0);
  assign w924[75] = |(datain[11:8] ^ 5);
  assign comp[924] = ~(|w924);
  wire [74-1:0] w925;
  assign w925[0] = |(datain[311:308] ^ 11);
  assign w925[1] = |(datain[307:304] ^ 10);
  assign w925[2] = |(datain[303:300] ^ 7);
  assign w925[3] = |(datain[299:296] ^ 1);
  assign w925[4] = |(datain[295:292] ^ 0);
  assign w925[5] = |(datain[291:288] ^ 0);
  assign w925[6] = |(datain[287:284] ^ 14);
  assign w925[7] = |(datain[283:280] ^ 12);
  assign w925[8] = |(datain[279:276] ^ 0);
  assign w925[9] = |(datain[275:272] ^ 12);
  assign w925[10] = |(datain[271:268] ^ 8);
  assign w925[11] = |(datain[267:264] ^ 0);
  assign w925[12] = |(datain[263:260] ^ 14);
  assign w925[13] = |(datain[259:256] ^ 14);
  assign w925[14] = |(datain[255:252] ^ 0);
  assign w925[15] = |(datain[251:248] ^ 7);
  assign w925[16] = |(datain[247:244] ^ 11);
  assign w925[17] = |(datain[243:240] ^ 14);
  assign w925[18] = |(datain[239:236] ^ 4);
  assign w925[19] = |(datain[235:232] ^ 12);
  assign w925[20] = |(datain[231:228] ^ 0);
  assign w925[21] = |(datain[227:224] ^ 0);
  assign w925[22] = |(datain[223:220] ^ 11);
  assign w925[23] = |(datain[219:216] ^ 15);
  assign w925[24] = |(datain[215:212] ^ 2);
  assign w925[25] = |(datain[211:208] ^ 11);
  assign w925[26] = |(datain[207:204] ^ 0);
  assign w925[27] = |(datain[203:200] ^ 1);
  assign w925[28] = |(datain[199:196] ^ 15);
  assign w925[29] = |(datain[195:192] ^ 12);
  assign w925[30] = |(datain[191:188] ^ 10);
  assign w925[31] = |(datain[187:184] ^ 5);
  assign w925[32] = |(datain[183:180] ^ 10);
  assign w925[33] = |(datain[179:176] ^ 5);
  assign w925[34] = |(datain[175:172] ^ 8);
  assign w925[35] = |(datain[171:168] ^ 12);
  assign w925[36] = |(datain[167:164] ^ 4);
  assign w925[37] = |(datain[163:160] ^ 4);
  assign w925[38] = |(datain[159:156] ^ 15);
  assign w925[39] = |(datain[155:152] ^ 14);
  assign w925[40] = |(datain[151:148] ^ 12);
  assign w925[41] = |(datain[147:144] ^ 7);
  assign w925[42] = |(datain[143:140] ^ 4);
  assign w925[43] = |(datain[139:136] ^ 4);
  assign w925[44] = |(datain[135:132] ^ 15);
  assign w925[45] = |(datain[131:128] ^ 12);
  assign w925[46] = |(datain[127:124] ^ 3);
  assign w925[47] = |(datain[123:120] ^ 1);
  assign w925[48] = |(datain[119:116] ^ 0);
  assign w925[49] = |(datain[115:112] ^ 1);
  assign w925[50] = |(datain[111:108] ^ 11);
  assign w925[51] = |(datain[107:104] ^ 4);
  assign w925[52] = |(datain[103:100] ^ 0);
  assign w925[53] = |(datain[99:96] ^ 4);
  assign w925[54] = |(datain[95:92] ^ 12);
  assign w925[55] = |(datain[91:88] ^ 13);
  assign w925[56] = |(datain[87:84] ^ 1);
  assign w925[57] = |(datain[83:80] ^ 10);
  assign w925[58] = |(datain[79:76] ^ 8);
  assign w925[59] = |(datain[75:72] ^ 1);
  assign w925[60] = |(datain[71:68] ^ 15);
  assign w925[61] = |(datain[67:64] ^ 10);
  assign w925[62] = |(datain[63:60] ^ 0);
  assign w925[63] = |(datain[59:56] ^ 4);
  assign w925[64] = |(datain[55:52] ^ 0);
  assign w925[65] = |(datain[51:48] ^ 9);
  assign w925[66] = |(datain[47:44] ^ 7);
  assign w925[67] = |(datain[43:40] ^ 5);
  assign w925[68] = |(datain[39:36] ^ 3);
  assign w925[69] = |(datain[35:32] ^ 9);
  assign w925[70] = |(datain[31:28] ^ 11);
  assign w925[71] = |(datain[27:24] ^ 4);
  assign w925[72] = |(datain[23:20] ^ 0);
  assign w925[73] = |(datain[19:16] ^ 6);
  assign comp[925] = ~(|w925);
  wire [76-1:0] w926;
  assign w926[0] = |(datain[311:308] ^ 1);
  assign w926[1] = |(datain[307:304] ^ 3);
  assign w926[2] = |(datain[303:300] ^ 7);
  assign w926[3] = |(datain[299:296] ^ 2);
  assign w926[4] = |(datain[295:292] ^ 1);
  assign w926[5] = |(datain[291:288] ^ 13);
  assign w926[6] = |(datain[287:284] ^ 11);
  assign w926[7] = |(datain[283:280] ^ 14);
  assign w926[8] = |(datain[279:276] ^ 11);
  assign w926[9] = |(datain[275:272] ^ 14);
  assign w926[10] = |(datain[271:268] ^ 8);
  assign w926[11] = |(datain[267:264] ^ 0);
  assign w926[12] = |(datain[263:260] ^ 11);
  assign w926[13] = |(datain[259:256] ^ 15);
  assign w926[14] = |(datain[255:252] ^ 11);
  assign w926[15] = |(datain[251:248] ^ 14);
  assign w926[16] = |(datain[247:244] ^ 7);
  assign w926[17] = |(datain[243:240] ^ 13);
  assign w926[18] = |(datain[239:236] ^ 11);
  assign w926[19] = |(datain[235:232] ^ 9);
  assign w926[20] = |(datain[231:228] ^ 2);
  assign w926[21] = |(datain[227:224] ^ 1);
  assign w926[22] = |(datain[223:220] ^ 0);
  assign w926[23] = |(datain[219:216] ^ 0);
  assign w926[24] = |(datain[215:212] ^ 15);
  assign w926[25] = |(datain[211:208] ^ 3);
  assign w926[26] = |(datain[207:204] ^ 10);
  assign w926[27] = |(datain[203:200] ^ 5);
  assign w926[28] = |(datain[199:196] ^ 5);
  assign w926[29] = |(datain[195:192] ^ 9);
  assign w926[30] = |(datain[191:188] ^ 8);
  assign w926[31] = |(datain[187:184] ^ 0);
  assign w926[32] = |(datain[183:180] ^ 3);
  assign w926[33] = |(datain[179:176] ^ 14);
  assign w926[34] = |(datain[175:172] ^ 11);
  assign w926[35] = |(datain[171:168] ^ 7);
  assign w926[36] = |(datain[167:164] ^ 7);
  assign w926[37] = |(datain[163:160] ^ 13);
  assign w926[38] = |(datain[159:156] ^ 0);
  assign w926[39] = |(datain[155:152] ^ 0);
  assign w926[40] = |(datain[151:148] ^ 7);
  assign w926[41] = |(datain[147:144] ^ 5);
  assign w926[42] = |(datain[143:140] ^ 0);
  assign w926[43] = |(datain[139:136] ^ 15);
  assign w926[44] = |(datain[135:132] ^ 11);
  assign w926[45] = |(datain[131:128] ^ 8);
  assign w926[46] = |(datain[127:124] ^ 0);
  assign w926[47] = |(datain[123:120] ^ 1);
  assign w926[48] = |(datain[119:116] ^ 0);
  assign w926[49] = |(datain[115:112] ^ 3);
  assign w926[50] = |(datain[111:108] ^ 11);
  assign w926[51] = |(datain[107:104] ^ 11);
  assign w926[52] = |(datain[103:100] ^ 0);
  assign w926[53] = |(datain[99:96] ^ 0);
  assign w926[54] = |(datain[95:92] ^ 7);
  assign w926[55] = |(datain[91:88] ^ 12);
  assign w926[56] = |(datain[87:84] ^ 12);
  assign w926[57] = |(datain[83:80] ^ 13);
  assign w926[58] = |(datain[79:76] ^ 1);
  assign w926[59] = |(datain[75:72] ^ 3);
  assign w926[60] = |(datain[71:68] ^ 7);
  assign w926[61] = |(datain[67:64] ^ 3);
  assign w926[62] = |(datain[63:60] ^ 0);
  assign w926[63] = |(datain[59:56] ^ 5);
  assign w926[64] = |(datain[55:52] ^ 11);
  assign w926[65] = |(datain[51:48] ^ 14);
  assign w926[66] = |(datain[47:44] ^ 8);
  assign w926[67] = |(datain[43:40] ^ 10);
  assign w926[68] = |(datain[39:36] ^ 7);
  assign w926[69] = |(datain[35:32] ^ 13);
  assign w926[70] = |(datain[31:28] ^ 14);
  assign w926[71] = |(datain[27:24] ^ 11);
  assign w926[72] = |(datain[23:20] ^ 5);
  assign w926[73] = |(datain[19:16] ^ 13);
  assign w926[74] = |(datain[15:12] ^ 15);
  assign w926[75] = |(datain[11:8] ^ 10);
  assign comp[926] = ~(|w926);
  wire [76-1:0] w927;
  assign w927[0] = |(datain[311:308] ^ 8);
  assign w927[1] = |(datain[307:304] ^ 3);
  assign w927[2] = |(datain[303:300] ^ 2);
  assign w927[3] = |(datain[299:296] ^ 14);
  assign w927[4] = |(datain[295:292] ^ 1);
  assign w927[5] = |(datain[291:288] ^ 3);
  assign w927[6] = |(datain[287:284] ^ 0);
  assign w927[7] = |(datain[283:280] ^ 4);
  assign w927[8] = |(datain[279:276] ^ 0);
  assign w927[9] = |(datain[275:272] ^ 8);
  assign w927[10] = |(datain[271:268] ^ 12);
  assign w927[11] = |(datain[267:264] ^ 13);
  assign w927[12] = |(datain[263:260] ^ 1);
  assign w927[13] = |(datain[259:256] ^ 2);
  assign w927[14] = |(datain[255:252] ^ 11);
  assign w927[15] = |(datain[251:248] ^ 1);
  assign w927[16] = |(datain[247:244] ^ 0);
  assign w927[17] = |(datain[243:240] ^ 6);
  assign w927[18] = |(datain[239:236] ^ 13);
  assign w927[19] = |(datain[235:232] ^ 3);
  assign w927[20] = |(datain[231:228] ^ 14);
  assign w927[21] = |(datain[227:224] ^ 0);
  assign w927[22] = |(datain[223:220] ^ 8);
  assign w927[23] = |(datain[219:216] ^ 14);
  assign w927[24] = |(datain[215:212] ^ 12);
  assign w927[25] = |(datain[211:208] ^ 0);
  assign w927[26] = |(datain[207:204] ^ 3);
  assign w927[27] = |(datain[203:200] ^ 3);
  assign w927[28] = |(datain[199:196] ^ 12);
  assign w927[29] = |(datain[195:192] ^ 0);
  assign w927[30] = |(datain[191:188] ^ 12);
  assign w927[31] = |(datain[187:184] ^ 13);
  assign w927[32] = |(datain[183:180] ^ 1);
  assign w927[33] = |(datain[179:176] ^ 3);
  assign w927[34] = |(datain[175:172] ^ 3);
  assign w927[35] = |(datain[171:168] ^ 2);
  assign w927[36] = |(datain[167:164] ^ 15);
  assign w927[37] = |(datain[163:160] ^ 6);
  assign w927[38] = |(datain[159:156] ^ 11);
  assign w927[39] = |(datain[155:152] ^ 9);
  assign w927[40] = |(datain[151:148] ^ 0);
  assign w927[41] = |(datain[147:144] ^ 4);
  assign w927[42] = |(datain[143:140] ^ 0);
  assign w927[43] = |(datain[139:136] ^ 0);
  assign w927[44] = |(datain[135:132] ^ 0);
  assign w927[45] = |(datain[131:128] ^ 10);
  assign w927[46] = |(datain[127:124] ^ 13);
  assign w927[47] = |(datain[123:120] ^ 2);
  assign w927[48] = |(datain[119:116] ^ 7);
  assign w927[49] = |(datain[115:112] ^ 8);
  assign w927[50] = |(datain[111:108] ^ 0);
  assign w927[51] = |(datain[107:104] ^ 5);
  assign w927[52] = |(datain[103:100] ^ 11);
  assign w927[53] = |(datain[99:96] ^ 9);
  assign w927[54] = |(datain[95:92] ^ 0);
  assign w927[55] = |(datain[91:88] ^ 4);
  assign w927[56] = |(datain[87:84] ^ 0);
  assign w927[57] = |(datain[83:80] ^ 0);
  assign w927[58] = |(datain[79:76] ^ 11);
  assign w927[59] = |(datain[75:72] ^ 6);
  assign w927[60] = |(datain[71:68] ^ 0);
  assign w927[61] = |(datain[67:64] ^ 0);
  assign w927[62] = |(datain[63:60] ^ 3);
  assign w927[63] = |(datain[59:56] ^ 3);
  assign w927[64] = |(datain[55:52] ^ 13);
  assign w927[65] = |(datain[51:48] ^ 11);
  assign w927[66] = |(datain[47:44] ^ 11);
  assign w927[67] = |(datain[43:40] ^ 8);
  assign w927[68] = |(datain[39:36] ^ 0);
  assign w927[69] = |(datain[35:32] ^ 7);
  assign w927[70] = |(datain[31:28] ^ 0);
  assign w927[71] = |(datain[27:24] ^ 2);
  assign w927[72] = |(datain[23:20] ^ 12);
  assign w927[73] = |(datain[19:16] ^ 13);
  assign w927[74] = |(datain[15:12] ^ 1);
  assign w927[75] = |(datain[11:8] ^ 3);
  assign comp[927] = ~(|w927);
  wire [46-1:0] w928;
  assign w928[0] = |(datain[311:308] ^ 8);
  assign w928[1] = |(datain[307:304] ^ 14);
  assign w928[2] = |(datain[303:300] ^ 13);
  assign w928[3] = |(datain[299:296] ^ 0);
  assign w928[4] = |(datain[295:292] ^ 11);
  assign w928[5] = |(datain[291:288] ^ 12);
  assign w928[6] = |(datain[287:284] ^ 0);
  assign w928[7] = |(datain[283:280] ^ 0);
  assign w928[8] = |(datain[279:276] ^ 7);
  assign w928[9] = |(datain[275:272] ^ 12);
  assign w928[10] = |(datain[271:268] ^ 1);
  assign w928[11] = |(datain[267:264] ^ 6);
  assign w928[12] = |(datain[263:260] ^ 0);
  assign w928[13] = |(datain[259:256] ^ 7);
  assign w928[14] = |(datain[255:252] ^ 11);
  assign w928[15] = |(datain[251:248] ^ 11);
  assign w928[16] = |(datain[247:244] ^ 0);
  assign w928[17] = |(datain[243:240] ^ 0);
  assign w928[18] = |(datain[239:236] ^ 7);
  assign w928[19] = |(datain[235:232] ^ 14);
  assign w928[20] = |(datain[231:228] ^ 11);
  assign w928[21] = |(datain[227:224] ^ 8);
  assign w928[22] = |(datain[223:220] ^ 0);
  assign w928[23] = |(datain[219:216] ^ 1);
  assign w928[24] = |(datain[215:212] ^ 0);
  assign w928[25] = |(datain[211:208] ^ 2);
  assign w928[26] = |(datain[207:204] ^ 11);
  assign w928[27] = |(datain[203:200] ^ 9);
  assign w928[28] = |(datain[199:196] ^ 0);
  assign w928[29] = |(datain[195:192] ^ 6);
  assign w928[30] = |(datain[191:188] ^ 2);
  assign w928[31] = |(datain[187:184] ^ 7);
  assign w928[32] = |(datain[183:180] ^ 11);
  assign w928[33] = |(datain[179:176] ^ 10);
  assign w928[34] = |(datain[175:172] ^ 0);
  assign w928[35] = |(datain[171:168] ^ 0);
  assign w928[36] = |(datain[167:164] ^ 0);
  assign w928[37] = |(datain[163:160] ^ 1);
  assign w928[38] = |(datain[159:156] ^ 12);
  assign w928[39] = |(datain[155:152] ^ 13);
  assign w928[40] = |(datain[151:148] ^ 1);
  assign w928[41] = |(datain[147:144] ^ 3);
  assign w928[42] = |(datain[143:140] ^ 15);
  assign w928[43] = |(datain[139:136] ^ 15);
  assign w928[44] = |(datain[135:132] ^ 14);
  assign w928[45] = |(datain[131:128] ^ 3);
  assign comp[928] = ~(|w928);
  wire [28-1:0] w929;
  assign w929[0] = |(datain[311:308] ^ 11);
  assign w929[1] = |(datain[307:304] ^ 9);
  assign w929[2] = |(datain[303:300] ^ 4);
  assign w929[3] = |(datain[299:296] ^ 14);
  assign w929[4] = |(datain[295:292] ^ 0);
  assign w929[5] = |(datain[291:288] ^ 1);
  assign w929[6] = |(datain[287:284] ^ 15);
  assign w929[7] = |(datain[283:280] ^ 12);
  assign w929[8] = |(datain[279:276] ^ 15);
  assign w929[9] = |(datain[275:272] ^ 3);
  assign w929[10] = |(datain[271:268] ^ 10);
  assign w929[11] = |(datain[267:264] ^ 4);
  assign w929[12] = |(datain[263:260] ^ 0);
  assign w929[13] = |(datain[259:256] ^ 6);
  assign w929[14] = |(datain[255:252] ^ 1);
  assign w929[15] = |(datain[251:248] ^ 15);
  assign w929[16] = |(datain[247:244] ^ 3);
  assign w929[17] = |(datain[243:240] ^ 1);
  assign w929[18] = |(datain[239:236] ^ 13);
  assign w929[19] = |(datain[235:232] ^ 2);
  assign w929[20] = |(datain[231:228] ^ 11);
  assign w929[21] = |(datain[227:224] ^ 8);
  assign w929[22] = |(datain[223:220] ^ 2);
  assign w929[23] = |(datain[219:216] ^ 1);
  assign w929[24] = |(datain[215:212] ^ 2);
  assign w929[25] = |(datain[211:208] ^ 5);
  assign w929[26] = |(datain[207:204] ^ 12);
  assign w929[27] = |(datain[203:200] ^ 13);
  assign comp[929] = ~(|w929);
  wire [30-1:0] w930;
  assign w930[0] = |(datain[311:308] ^ 3);
  assign w930[1] = |(datain[307:304] ^ 13);
  assign w930[2] = |(datain[303:300] ^ 0);
  assign w930[3] = |(datain[299:296] ^ 0);
  assign w930[4] = |(datain[295:292] ^ 4);
  assign w930[5] = |(datain[291:288] ^ 11);
  assign w930[6] = |(datain[287:284] ^ 7);
  assign w930[7] = |(datain[283:280] ^ 5);
  assign w930[8] = |(datain[279:276] ^ 1);
  assign w930[9] = |(datain[275:272] ^ 0);
  assign w930[10] = |(datain[271:268] ^ 5);
  assign w930[11] = |(datain[267:264] ^ 6);
  assign w930[12] = |(datain[263:260] ^ 8);
  assign w930[13] = |(datain[259:256] ^ 9);
  assign w930[14] = |(datain[255:252] ^ 13);
  assign w930[15] = |(datain[251:248] ^ 6);
  assign w930[16] = |(datain[247:244] ^ 4);
  assign w930[17] = |(datain[243:240] ^ 6);
  assign w930[18] = |(datain[239:236] ^ 8);
  assign w930[19] = |(datain[235:232] ^ 0);
  assign w930[20] = |(datain[231:228] ^ 3);
  assign w930[21] = |(datain[227:224] ^ 12);
  assign w930[22] = |(datain[223:220] ^ 0);
  assign w930[23] = |(datain[219:216] ^ 0);
  assign w930[24] = |(datain[215:212] ^ 7);
  assign w930[25] = |(datain[211:208] ^ 5);
  assign w930[26] = |(datain[207:204] ^ 15);
  assign w930[27] = |(datain[203:200] ^ 10);
  assign w930[28] = |(datain[199:196] ^ 8);
  assign w930[29] = |(datain[195:192] ^ 0);
  assign comp[930] = ~(|w930);
  wire [46-1:0] w931;
  assign w931[0] = |(datain[311:308] ^ 3);
  assign w931[1] = |(datain[307:304] ^ 13);
  assign w931[2] = |(datain[303:300] ^ 0);
  assign w931[3] = |(datain[299:296] ^ 0);
  assign w931[4] = |(datain[295:292] ^ 4);
  assign w931[5] = |(datain[291:288] ^ 11);
  assign w931[6] = |(datain[287:284] ^ 7);
  assign w931[7] = |(datain[283:280] ^ 5);
  assign w931[8] = |(datain[279:276] ^ 1);
  assign w931[9] = |(datain[275:272] ^ 0);
  assign w931[10] = |(datain[271:268] ^ 5);
  assign w931[11] = |(datain[267:264] ^ 6);
  assign w931[12] = |(datain[263:260] ^ 8);
  assign w931[13] = |(datain[259:256] ^ 9);
  assign w931[14] = |(datain[255:252] ^ 13);
  assign w931[15] = |(datain[251:248] ^ 6);
  assign w931[16] = |(datain[247:244] ^ 4);
  assign w931[17] = |(datain[243:240] ^ 6);
  assign w931[18] = |(datain[239:236] ^ 8);
  assign w931[19] = |(datain[235:232] ^ 0);
  assign w931[20] = |(datain[231:228] ^ 3);
  assign w931[21] = |(datain[227:224] ^ 12);
  assign w931[22] = |(datain[223:220] ^ 0);
  assign w931[23] = |(datain[219:216] ^ 0);
  assign w931[24] = |(datain[215:212] ^ 7);
  assign w931[25] = |(datain[211:208] ^ 5);
  assign w931[26] = |(datain[207:204] ^ 15);
  assign w931[27] = |(datain[203:200] ^ 10);
  assign w931[28] = |(datain[199:196] ^ 8);
  assign w931[29] = |(datain[195:192] ^ 0);
  assign w931[30] = |(datain[191:188] ^ 7);
  assign w931[31] = |(datain[187:184] ^ 12);
  assign w931[32] = |(datain[183:180] ^ 15);
  assign w931[33] = |(datain[179:176] ^ 15);
  assign w931[34] = |(datain[175:172] ^ 4);
  assign w931[35] = |(datain[171:168] ^ 5);
  assign w931[36] = |(datain[167:164] ^ 7);
  assign w931[37] = |(datain[163:160] ^ 4);
  assign w931[38] = |(datain[159:156] ^ 0);
  assign w931[39] = |(datain[155:152] ^ 7);
  assign w931[40] = |(datain[151:148] ^ 5);
  assign w931[41] = |(datain[147:144] ^ 14);
  assign w931[42] = |(datain[143:140] ^ 9);
  assign w931[43] = |(datain[139:136] ^ 13);
  assign w931[44] = |(datain[135:132] ^ 14);
  assign w931[45] = |(datain[131:128] ^ 10);
  assign comp[931] = ~(|w931);
  wire [74-1:0] w932;
  assign w932[0] = |(datain[311:308] ^ 11);
  assign w932[1] = |(datain[307:304] ^ 1);
  assign w932[2] = |(datain[303:300] ^ 0);
  assign w932[3] = |(datain[299:296] ^ 6);
  assign w932[4] = |(datain[295:292] ^ 13);
  assign w932[5] = |(datain[291:288] ^ 3);
  assign w932[6] = |(datain[287:284] ^ 14);
  assign w932[7] = |(datain[283:280] ^ 0);
  assign w932[8] = |(datain[279:276] ^ 2);
  assign w932[9] = |(datain[275:272] ^ 14);
  assign w932[10] = |(datain[271:268] ^ 10);
  assign w932[11] = |(datain[267:264] ^ 3);
  assign w932[12] = |(datain[263:260] ^ 4);
  assign w932[13] = |(datain[259:256] ^ 4);
  assign w932[14] = |(datain[255:252] ^ 0);
  assign w932[15] = |(datain[251:248] ^ 0);
  assign w932[16] = |(datain[247:244] ^ 8);
  assign w932[17] = |(datain[243:240] ^ 14);
  assign w932[18] = |(datain[239:236] ^ 12);
  assign w932[19] = |(datain[235:232] ^ 0);
  assign w932[20] = |(datain[231:228] ^ 0);
  assign w932[21] = |(datain[227:224] ^ 5);
  assign w932[22] = |(datain[223:220] ^ 8);
  assign w932[23] = |(datain[219:216] ^ 0);
  assign w932[24] = |(datain[215:212] ^ 0);
  assign w932[25] = |(datain[211:208] ^ 0);
  assign w932[26] = |(datain[207:204] ^ 2);
  assign w932[27] = |(datain[203:200] ^ 14);
  assign w932[28] = |(datain[199:196] ^ 10);
  assign w932[29] = |(datain[195:192] ^ 3);
  assign w932[30] = |(datain[191:188] ^ 4);
  assign w932[31] = |(datain[187:184] ^ 2);
  assign w932[32] = |(datain[183:180] ^ 0);
  assign w932[33] = |(datain[179:176] ^ 0);
  assign w932[34] = |(datain[175:172] ^ 3);
  assign w932[35] = |(datain[171:168] ^ 3);
  assign w932[36] = |(datain[167:164] ^ 13);
  assign w932[37] = |(datain[163:160] ^ 11);
  assign w932[38] = |(datain[159:156] ^ 11);
  assign w932[39] = |(datain[155:152] ^ 8);
  assign w932[40] = |(datain[151:148] ^ 0);
  assign w932[41] = |(datain[147:144] ^ 6);
  assign w932[42] = |(datain[143:140] ^ 0);
  assign w932[43] = |(datain[139:136] ^ 2);
  assign w932[44] = |(datain[135:132] ^ 2);
  assign w932[45] = |(datain[131:128] ^ 14);
  assign w932[46] = |(datain[127:124] ^ 8);
  assign w932[47] = |(datain[123:120] ^ 0);
  assign w932[48] = |(datain[119:116] ^ 3);
  assign w932[49] = |(datain[115:112] ^ 14);
  assign w932[50] = |(datain[111:108] ^ 3);
  assign w932[51] = |(datain[107:104] ^ 14);
  assign w932[52] = |(datain[103:100] ^ 0);
  assign w932[53] = |(datain[99:96] ^ 0);
  assign w932[54] = |(datain[95:92] ^ 0);
  assign w932[55] = |(datain[91:88] ^ 0);
  assign w932[56] = |(datain[87:84] ^ 7);
  assign w932[57] = |(datain[83:80] ^ 4);
  assign w932[58] = |(datain[79:76] ^ 0);
  assign w932[59] = |(datain[75:72] ^ 10);
  assign w932[60] = |(datain[71:68] ^ 11);
  assign w932[61] = |(datain[67:64] ^ 9);
  assign w932[62] = |(datain[63:60] ^ 0);
  assign w932[63] = |(datain[59:56] ^ 8);
  assign w932[64] = |(datain[55:52] ^ 0);
  assign w932[65] = |(datain[51:48] ^ 0);
  assign w932[66] = |(datain[47:44] ^ 11);
  assign w932[67] = |(datain[43:40] ^ 10);
  assign w932[68] = |(datain[39:36] ^ 8);
  assign w932[69] = |(datain[35:32] ^ 0);
  assign w932[70] = |(datain[31:28] ^ 0);
  assign w932[71] = |(datain[27:24] ^ 0);
  assign w932[72] = |(datain[23:20] ^ 12);
  assign w932[73] = |(datain[19:16] ^ 13);
  assign comp[932] = ~(|w932);
  wire [74-1:0] w933;
  assign w933[0] = |(datain[311:308] ^ 12);
  assign w933[1] = |(datain[307:304] ^ 0);
  assign w933[2] = |(datain[303:300] ^ 0);
  assign w933[3] = |(datain[299:296] ^ 7);
  assign w933[4] = |(datain[295:292] ^ 3);
  assign w933[5] = |(datain[291:288] ^ 3);
  assign w933[6] = |(datain[287:284] ^ 12);
  assign w933[7] = |(datain[283:280] ^ 0);
  assign w933[8] = |(datain[279:276] ^ 8);
  assign w933[9] = |(datain[275:272] ^ 14);
  assign w933[10] = |(datain[271:268] ^ 13);
  assign w933[11] = |(datain[267:264] ^ 8);
  assign w933[12] = |(datain[263:260] ^ 8);
  assign w933[13] = |(datain[259:256] ^ 14);
  assign w933[14] = |(datain[255:252] ^ 13);
  assign w933[15] = |(datain[251:248] ^ 0);
  assign w933[16] = |(datain[247:244] ^ 11);
  assign w933[17] = |(datain[243:240] ^ 12);
  assign w933[18] = |(datain[239:236] ^ 0);
  assign w933[19] = |(datain[235:232] ^ 0);
  assign w933[20] = |(datain[231:228] ^ 7);
  assign w933[21] = |(datain[227:224] ^ 12);
  assign w933[22] = |(datain[223:220] ^ 2);
  assign w933[23] = |(datain[219:216] ^ 14);
  assign w933[24] = |(datain[215:212] ^ 8);
  assign w933[25] = |(datain[211:208] ^ 8);
  assign w933[26] = |(datain[207:204] ^ 1);
  assign w933[27] = |(datain[203:200] ^ 6);
  assign w933[28] = |(datain[199:196] ^ 1);
  assign w933[29] = |(datain[195:192] ^ 14);
  assign w933[30] = |(datain[191:188] ^ 0);
  assign w933[31] = |(datain[187:184] ^ 0);
  assign w933[32] = |(datain[183:180] ^ 15);
  assign w933[33] = |(datain[179:176] ^ 10);
  assign w933[34] = |(datain[175:172] ^ 10);
  assign w933[35] = |(datain[171:168] ^ 1);
  assign w933[36] = |(datain[167:164] ^ 4);
  assign w933[37] = |(datain[163:160] ^ 12);
  assign w933[38] = |(datain[159:156] ^ 0);
  assign w933[39] = |(datain[155:152] ^ 0);
  assign w933[40] = |(datain[151:148] ^ 8);
  assign w933[41] = |(datain[147:144] ^ 11);
  assign w933[42] = |(datain[143:140] ^ 1);
  assign w933[43] = |(datain[139:136] ^ 14);
  assign w933[44] = |(datain[135:132] ^ 4);
  assign w933[45] = |(datain[131:128] ^ 14);
  assign w933[46] = |(datain[127:124] ^ 0);
  assign w933[47] = |(datain[123:120] ^ 0);
  assign w933[48] = |(datain[119:116] ^ 2);
  assign w933[49] = |(datain[115:112] ^ 14);
  assign w933[50] = |(datain[111:108] ^ 10);
  assign w933[51] = |(datain[107:104] ^ 3);
  assign w933[52] = |(datain[103:100] ^ 2);
  assign w933[53] = |(datain[99:96] ^ 4);
  assign w933[54] = |(datain[95:92] ^ 0);
  assign w933[55] = |(datain[91:88] ^ 0);
  assign w933[56] = |(datain[87:84] ^ 2);
  assign w933[57] = |(datain[83:80] ^ 14);
  assign w933[58] = |(datain[79:76] ^ 8);
  assign w933[59] = |(datain[75:72] ^ 9);
  assign w933[60] = |(datain[71:68] ^ 1);
  assign w933[61] = |(datain[67:64] ^ 14);
  assign w933[62] = |(datain[63:60] ^ 2);
  assign w933[63] = |(datain[59:56] ^ 6);
  assign w933[64] = |(datain[55:52] ^ 0);
  assign w933[65] = |(datain[51:48] ^ 0);
  assign w933[66] = |(datain[47:44] ^ 15);
  assign w933[67] = |(datain[43:40] ^ 11);
  assign w933[68] = |(datain[39:36] ^ 10);
  assign w933[69] = |(datain[35:32] ^ 1);
  assign w933[70] = |(datain[31:28] ^ 1);
  assign w933[71] = |(datain[27:24] ^ 3);
  assign w933[72] = |(datain[23:20] ^ 0);
  assign w933[73] = |(datain[19:16] ^ 4);
  assign comp[933] = ~(|w933);
  wire [76-1:0] w934;
  assign w934[0] = |(datain[311:308] ^ 9);
  assign w934[1] = |(datain[307:304] ^ 3);
  assign w934[2] = |(datain[303:300] ^ 11);
  assign w934[3] = |(datain[299:296] ^ 10);
  assign w934[4] = |(datain[295:292] ^ 8);
  assign w934[5] = |(datain[291:288] ^ 0);
  assign w934[6] = |(datain[287:284] ^ 0);
  assign w934[7] = |(datain[283:280] ^ 0);
  assign w934[8] = |(datain[279:276] ^ 12);
  assign w934[9] = |(datain[275:272] ^ 13);
  assign w934[10] = |(datain[271:268] ^ 1);
  assign w934[11] = |(datain[267:264] ^ 3);
  assign w934[12] = |(datain[263:260] ^ 12);
  assign w934[13] = |(datain[259:256] ^ 7);
  assign w934[14] = |(datain[255:252] ^ 4);
  assign w934[15] = |(datain[251:248] ^ 7);
  assign w934[16] = |(datain[247:244] ^ 15);
  assign w934[17] = |(datain[243:240] ^ 14);
  assign w934[18] = |(datain[239:236] ^ 5);
  assign w934[19] = |(datain[235:232] ^ 5);
  assign w934[20] = |(datain[231:228] ^ 10);
  assign w934[21] = |(datain[227:224] ^ 10);
  assign w934[22] = |(datain[223:220] ^ 9);
  assign w934[23] = |(datain[219:216] ^ 6);
  assign w934[24] = |(datain[215:212] ^ 3);
  assign w934[25] = |(datain[211:208] ^ 8);
  assign w934[26] = |(datain[207:204] ^ 1);
  assign w934[27] = |(datain[203:200] ^ 15);
  assign w934[28] = |(datain[199:196] ^ 11);
  assign w934[29] = |(datain[195:192] ^ 3);
  assign w934[30] = |(datain[191:188] ^ 0);
  assign w934[31] = |(datain[187:184] ^ 2);
  assign w934[32] = |(datain[183:180] ^ 7);
  assign w934[33] = |(datain[179:176] ^ 5);
  assign w934[34] = |(datain[175:172] ^ 14);
  assign w934[35] = |(datain[171:168] ^ 14);
  assign w934[36] = |(datain[167:164] ^ 12);
  assign w934[37] = |(datain[163:160] ^ 3);
  assign w934[38] = |(datain[159:156] ^ 0);
  assign w934[39] = |(datain[155:152] ^ 14);
  assign w934[40] = |(datain[151:148] ^ 1);
  assign w934[41] = |(datain[147:144] ^ 15);
  assign w934[42] = |(datain[143:140] ^ 8);
  assign w934[43] = |(datain[139:136] ^ 7);
  assign w934[44] = |(datain[135:132] ^ 13);
  assign w934[45] = |(datain[131:128] ^ 14);
  assign w934[46] = |(datain[127:124] ^ 15);
  assign w934[47] = |(datain[123:120] ^ 15);
  assign w934[48] = |(datain[119:116] ^ 0);
  assign w934[49] = |(datain[115:112] ^ 14);
  assign w934[50] = |(datain[111:108] ^ 1);
  assign w934[51] = |(datain[107:104] ^ 3);
  assign w934[52] = |(datain[103:100] ^ 0);
  assign w934[53] = |(datain[99:96] ^ 4);
  assign w934[54] = |(datain[95:92] ^ 12);
  assign w934[55] = |(datain[91:88] ^ 13);
  assign w934[56] = |(datain[87:84] ^ 1);
  assign w934[57] = |(datain[83:80] ^ 2);
  assign w934[58] = |(datain[79:76] ^ 11);
  assign w934[59] = |(datain[75:72] ^ 1);
  assign w934[60] = |(datain[71:68] ^ 7);
  assign w934[61] = |(datain[67:64] ^ 6);
  assign w934[62] = |(datain[63:60] ^ 13);
  assign w934[63] = |(datain[59:56] ^ 3);
  assign w934[64] = |(datain[55:52] ^ 12);
  assign w934[65] = |(datain[51:48] ^ 0);
  assign w934[66] = |(datain[47:44] ^ 8);
  assign w934[67] = |(datain[43:40] ^ 14);
  assign w934[68] = |(datain[39:36] ^ 12);
  assign w934[69] = |(datain[35:32] ^ 0);
  assign w934[70] = |(datain[31:28] ^ 3);
  assign w934[71] = |(datain[27:24] ^ 3);
  assign w934[72] = |(datain[23:20] ^ 15);
  assign w934[73] = |(datain[19:16] ^ 15);
  assign w934[74] = |(datain[15:12] ^ 15);
  assign w934[75] = |(datain[11:8] ^ 3);
  assign comp[934] = ~(|w934);
  wire [76-1:0] w935;
  assign w935[0] = |(datain[311:308] ^ 7);
  assign w935[1] = |(datain[307:304] ^ 12);
  assign w935[2] = |(datain[303:300] ^ 15);
  assign w935[3] = |(datain[299:296] ^ 11);
  assign w935[4] = |(datain[295:292] ^ 15);
  assign w935[5] = |(datain[291:288] ^ 12);
  assign w935[6] = |(datain[287:284] ^ 1);
  assign w935[7] = |(datain[283:280] ^ 6);
  assign w935[8] = |(datain[279:276] ^ 1);
  assign w935[9] = |(datain[275:272] ^ 15);
  assign w935[10] = |(datain[271:268] ^ 12);
  assign w935[11] = |(datain[267:264] ^ 13);
  assign w935[12] = |(datain[263:260] ^ 1);
  assign w935[13] = |(datain[259:256] ^ 2);
  assign w935[14] = |(datain[255:252] ^ 2);
  assign w935[15] = |(datain[251:248] ^ 13);
  assign w935[16] = |(datain[247:244] ^ 0);
  assign w935[17] = |(datain[243:240] ^ 11);
  assign w935[18] = |(datain[239:236] ^ 0);
  assign w935[19] = |(datain[235:232] ^ 0);
  assign w935[20] = |(datain[231:228] ^ 10);
  assign w935[21] = |(datain[227:224] ^ 3);
  assign w935[22] = |(datain[223:220] ^ 1);
  assign w935[23] = |(datain[219:216] ^ 3);
  assign w935[24] = |(datain[215:212] ^ 0);
  assign w935[25] = |(datain[211:208] ^ 4);
  assign w935[26] = |(datain[207:204] ^ 11);
  assign w935[27] = |(datain[203:200] ^ 1);
  assign w935[28] = |(datain[199:196] ^ 0);
  assign w935[29] = |(datain[195:192] ^ 6);
  assign w935[30] = |(datain[191:188] ^ 13);
  assign w935[31] = |(datain[187:184] ^ 3);
  assign w935[32] = |(datain[183:180] ^ 14);
  assign w935[33] = |(datain[179:176] ^ 0);
  assign w935[34] = |(datain[175:172] ^ 8);
  assign w935[35] = |(datain[171:168] ^ 14);
  assign w935[36] = |(datain[167:164] ^ 12);
  assign w935[37] = |(datain[163:160] ^ 0);
  assign w935[38] = |(datain[159:156] ^ 11);
  assign w935[39] = |(datain[155:152] ^ 14);
  assign w935[40] = |(datain[151:148] ^ 0);
  assign w935[41] = |(datain[147:144] ^ 0);
  assign w935[42] = |(datain[143:140] ^ 7);
  assign w935[43] = |(datain[139:136] ^ 12);
  assign w935[44] = |(datain[135:132] ^ 3);
  assign w935[45] = |(datain[131:128] ^ 3);
  assign w935[46] = |(datain[127:124] ^ 15);
  assign w935[47] = |(datain[123:120] ^ 15);
  assign w935[48] = |(datain[119:116] ^ 11);
  assign w935[49] = |(datain[115:112] ^ 9);
  assign w935[50] = |(datain[111:108] ^ 0);
  assign w935[51] = |(datain[107:104] ^ 0);
  assign w935[52] = |(datain[103:100] ^ 0);
  assign w935[53] = |(datain[99:96] ^ 1);
  assign w935[54] = |(datain[95:92] ^ 15);
  assign w935[55] = |(datain[91:88] ^ 3);
  assign w935[56] = |(datain[87:84] ^ 10);
  assign w935[57] = |(datain[83:80] ^ 5);
  assign w935[58] = |(datain[79:76] ^ 11);
  assign w935[59] = |(datain[75:72] ^ 8);
  assign w935[60] = |(datain[71:68] ^ 0);
  assign w935[61] = |(datain[67:64] ^ 8);
  assign w935[62] = |(datain[63:60] ^ 0);
  assign w935[63] = |(datain[59:56] ^ 2);
  assign w935[64] = |(datain[55:52] ^ 11);
  assign w935[65] = |(datain[51:48] ^ 11);
  assign w935[66] = |(datain[47:44] ^ 0);
  assign w935[67] = |(datain[43:40] ^ 0);
  assign w935[68] = |(datain[39:36] ^ 0);
  assign w935[69] = |(datain[35:32] ^ 2);
  assign w935[70] = |(datain[31:28] ^ 2);
  assign w935[71] = |(datain[27:24] ^ 6);
  assign w935[72] = |(datain[23:20] ^ 8);
  assign w935[73] = |(datain[19:16] ^ 0);
  assign w935[74] = |(datain[15:12] ^ 3);
  assign w935[75] = |(datain[11:8] ^ 14);
  assign comp[935] = ~(|w935);
  wire [54-1:0] w936;
  assign w936[0] = |(datain[311:308] ^ 11);
  assign w936[1] = |(datain[307:304] ^ 8);
  assign w936[2] = |(datain[303:300] ^ 0);
  assign w936[3] = |(datain[299:296] ^ 0);
  assign w936[4] = |(datain[295:292] ^ 0);
  assign w936[5] = |(datain[291:288] ^ 0);
  assign w936[6] = |(datain[287:284] ^ 11);
  assign w936[7] = |(datain[283:280] ^ 12);
  assign w936[8] = |(datain[279:276] ^ 0);
  assign w936[9] = |(datain[275:272] ^ 0);
  assign w936[10] = |(datain[271:268] ^ 7);
  assign w936[11] = |(datain[267:264] ^ 12);
  assign w936[12] = |(datain[263:260] ^ 8);
  assign w936[13] = |(datain[259:256] ^ 14);
  assign w936[14] = |(datain[255:252] ^ 13);
  assign w936[15] = |(datain[251:248] ^ 0);
  assign w936[16] = |(datain[247:244] ^ 1);
  assign w936[17] = |(datain[243:240] ^ 6);
  assign w936[18] = |(datain[239:236] ^ 0);
  assign w936[19] = |(datain[235:232] ^ 7);
  assign w936[20] = |(datain[231:228] ^ 11);
  assign w936[21] = |(datain[227:224] ^ 8);
  assign w936[22] = |(datain[223:220] ^ 0);
  assign w936[23] = |(datain[219:216] ^ 3);
  assign w936[24] = |(datain[215:212] ^ 0);
  assign w936[25] = |(datain[211:208] ^ 2);
  assign w936[26] = |(datain[207:204] ^ 11);
  assign w936[27] = |(datain[203:200] ^ 11);
  assign w936[28] = |(datain[199:196] ^ 0);
  assign w936[29] = |(datain[195:192] ^ 0);
  assign w936[30] = |(datain[191:188] ^ 7);
  assign w936[31] = |(datain[187:184] ^ 14);
  assign w936[32] = |(datain[183:180] ^ 11);
  assign w936[33] = |(datain[179:176] ^ 9);
  assign w936[34] = |(datain[175:172] ^ 0);
  assign w936[35] = |(datain[171:168] ^ 2);
  assign w936[36] = |(datain[167:164] ^ 0);
  assign w936[37] = |(datain[163:160] ^ 0);
  assign w936[38] = |(datain[159:156] ^ 11);
  assign w936[39] = |(datain[155:152] ^ 10);
  assign w936[40] = |(datain[151:148] ^ 0);
  assign w936[41] = |(datain[147:144] ^ 0);
  assign w936[42] = |(datain[143:140] ^ 0);
  assign w936[43] = |(datain[139:136] ^ 0);
  assign w936[44] = |(datain[135:132] ^ 12);
  assign w936[45] = |(datain[131:128] ^ 13);
  assign w936[46] = |(datain[127:124] ^ 1);
  assign w936[47] = |(datain[123:120] ^ 3);
  assign w936[48] = |(datain[119:116] ^ 14);
  assign w936[49] = |(datain[115:112] ^ 9);
  assign w936[50] = |(datain[111:108] ^ 9);
  assign w936[51] = |(datain[107:104] ^ 6);
  assign w936[52] = |(datain[103:100] ^ 0);
  assign w936[53] = |(datain[99:96] ^ 1);
  assign comp[936] = ~(|w936);
  wire [76-1:0] w937;
  assign w937[0] = |(datain[311:308] ^ 0);
  assign w937[1] = |(datain[307:304] ^ 2);
  assign w937[2] = |(datain[303:300] ^ 11);
  assign w937[3] = |(datain[299:296] ^ 9);
  assign w937[4] = |(datain[295:292] ^ 0);
  assign w937[5] = |(datain[291:288] ^ 7);
  assign w937[6] = |(datain[287:284] ^ 0);
  assign w937[7] = |(datain[283:280] ^ 0);
  assign w937[8] = |(datain[279:276] ^ 8);
  assign w937[9] = |(datain[275:272] ^ 9);
  assign w937[10] = |(datain[271:268] ^ 0);
  assign w937[11] = |(datain[267:264] ^ 14);
  assign w937[12] = |(datain[263:260] ^ 9);
  assign w937[13] = |(datain[259:256] ^ 3);
  assign w937[14] = |(datain[255:252] ^ 0);
  assign w937[15] = |(datain[251:248] ^ 1);
  assign w937[16] = |(datain[247:244] ^ 11);
  assign w937[17] = |(datain[243:240] ^ 8);
  assign w937[18] = |(datain[239:236] ^ 0);
  assign w937[19] = |(datain[235:232] ^ 1);
  assign w937[20] = |(datain[231:228] ^ 0);
  assign w937[21] = |(datain[227:224] ^ 3);
  assign w937[22] = |(datain[223:220] ^ 11);
  assign w937[23] = |(datain[219:216] ^ 10);
  assign w937[24] = |(datain[215:212] ^ 8);
  assign w937[25] = |(datain[211:208] ^ 0);
  assign w937[26] = |(datain[207:204] ^ 0);
  assign w937[27] = |(datain[203:200] ^ 0);
  assign w937[28] = |(datain[199:196] ^ 12);
  assign w937[29] = |(datain[195:192] ^ 13);
  assign w937[30] = |(datain[191:188] ^ 1);
  assign w937[31] = |(datain[187:184] ^ 3);
  assign w937[32] = |(datain[183:180] ^ 7);
  assign w937[33] = |(datain[179:176] ^ 2);
  assign w937[34] = |(datain[175:172] ^ 10);
  assign w937[35] = |(datain[171:168] ^ 10);
  assign w937[36] = |(datain[167:164] ^ 11);
  assign w937[37] = |(datain[163:160] ^ 14);
  assign w937[38] = |(datain[159:156] ^ 9);
  assign w937[39] = |(datain[155:152] ^ 11);
  assign w937[40] = |(datain[151:148] ^ 0);
  assign w937[41] = |(datain[147:144] ^ 3);
  assign w937[42] = |(datain[143:140] ^ 11);
  assign w937[43] = |(datain[139:136] ^ 15);
  assign w937[44] = |(datain[135:132] ^ 9);
  assign w937[45] = |(datain[131:128] ^ 11);
  assign w937[46] = |(datain[127:124] ^ 0);
  assign w937[47] = |(datain[123:120] ^ 1);
  assign w937[48] = |(datain[119:116] ^ 11);
  assign w937[49] = |(datain[115:112] ^ 9);
  assign w937[50] = |(datain[111:108] ^ 6);
  assign w937[51] = |(datain[107:104] ^ 9);
  assign w937[52] = |(datain[103:100] ^ 0);
  assign w937[53] = |(datain[99:96] ^ 0);
  assign w937[54] = |(datain[95:92] ^ 15);
  assign w937[55] = |(datain[91:88] ^ 3);
  assign w937[56] = |(datain[87:84] ^ 10);
  assign w937[57] = |(datain[83:80] ^ 4);
  assign w937[58] = |(datain[79:76] ^ 11);
  assign w937[59] = |(datain[75:72] ^ 8);
  assign w937[60] = |(datain[71:68] ^ 0);
  assign w937[61] = |(datain[67:64] ^ 1);
  assign w937[62] = |(datain[63:60] ^ 0);
  assign w937[63] = |(datain[59:56] ^ 3);
  assign w937[64] = |(datain[55:52] ^ 3);
  assign w937[65] = |(datain[51:48] ^ 3);
  assign w937[66] = |(datain[47:44] ^ 13);
  assign w937[67] = |(datain[43:40] ^ 11);
  assign w937[68] = |(datain[39:36] ^ 15);
  assign w937[69] = |(datain[35:32] ^ 14);
  assign w937[70] = |(datain[31:28] ^ 12);
  assign w937[71] = |(datain[27:24] ^ 1);
  assign w937[72] = |(datain[23:20] ^ 12);
  assign w937[73] = |(datain[19:16] ^ 13);
  assign w937[74] = |(datain[15:12] ^ 1);
  assign w937[75] = |(datain[11:8] ^ 3);
  assign comp[937] = ~(|w937);
  wire [74-1:0] w938;
  assign w938[0] = |(datain[311:308] ^ 4);
  assign w938[1] = |(datain[307:304] ^ 12);
  assign w938[2] = |(datain[303:300] ^ 0);
  assign w938[3] = |(datain[299:296] ^ 0);
  assign w938[4] = |(datain[295:292] ^ 8);
  assign w938[5] = |(datain[291:288] ^ 15);
  assign w938[6] = |(datain[287:284] ^ 0);
  assign w938[7] = |(datain[283:280] ^ 6);
  assign w938[8] = |(datain[279:276] ^ 4);
  assign w938[9] = |(datain[275:272] ^ 14);
  assign w938[10] = |(datain[271:268] ^ 0);
  assign w938[11] = |(datain[267:264] ^ 0);
  assign w938[12] = |(datain[263:260] ^ 12);
  assign w938[13] = |(datain[259:256] ^ 7);
  assign w938[14] = |(datain[255:252] ^ 0);
  assign w938[15] = |(datain[251:248] ^ 6);
  assign w938[16] = |(datain[247:244] ^ 6);
  assign w938[17] = |(datain[243:240] ^ 0);
  assign w938[18] = |(datain[239:236] ^ 0);
  assign w938[19] = |(datain[235:232] ^ 0);
  assign w938[20] = |(datain[231:228] ^ 1);
  assign w938[21] = |(datain[227:224] ^ 11);
  assign w938[22] = |(datain[223:220] ^ 0);
  assign w938[23] = |(datain[219:216] ^ 1);
  assign w938[24] = |(datain[215:212] ^ 8);
  assign w938[25] = |(datain[211:208] ^ 12);
  assign w938[26] = |(datain[207:204] ^ 0);
  assign w938[27] = |(datain[203:200] ^ 6);
  assign w938[28] = |(datain[199:196] ^ 6);
  assign w938[29] = |(datain[195:192] ^ 2);
  assign w938[30] = |(datain[191:188] ^ 0);
  assign w938[31] = |(datain[187:184] ^ 0);
  assign w938[32] = |(datain[183:180] ^ 0);
  assign w938[33] = |(datain[179:176] ^ 14);
  assign w938[34] = |(datain[175:172] ^ 0);
  assign w938[35] = |(datain[171:168] ^ 7);
  assign w938[36] = |(datain[167:164] ^ 11);
  assign w938[37] = |(datain[163:160] ^ 11);
  assign w938[38] = |(datain[159:156] ^ 0);
  assign w938[39] = |(datain[155:152] ^ 0);
  assign w938[40] = |(datain[151:148] ^ 0);
  assign w938[41] = |(datain[147:144] ^ 2);
  assign w938[42] = |(datain[143:140] ^ 11);
  assign w938[43] = |(datain[139:136] ^ 9);
  assign w938[44] = |(datain[135:132] ^ 0);
  assign w938[45] = |(datain[131:128] ^ 8);
  assign w938[46] = |(datain[127:124] ^ 0);
  assign w938[47] = |(datain[123:120] ^ 0);
  assign w938[48] = |(datain[119:116] ^ 3);
  assign w938[49] = |(datain[115:112] ^ 2);
  assign w938[50] = |(datain[111:108] ^ 15);
  assign w938[51] = |(datain[107:104] ^ 6);
  assign w938[52] = |(datain[103:100] ^ 14);
  assign w938[53] = |(datain[99:96] ^ 8);
  assign w938[54] = |(datain[95:92] ^ 5);
  assign w938[55] = |(datain[91:88] ^ 15);
  assign w938[56] = |(datain[87:84] ^ 0);
  assign w938[57] = |(datain[83:80] ^ 0);
  assign w938[58] = |(datain[79:76] ^ 11);
  assign w938[59] = |(datain[75:72] ^ 4);
  assign w938[60] = |(datain[71:68] ^ 0);
  assign w938[61] = |(datain[67:64] ^ 4);
  assign w938[62] = |(datain[63:60] ^ 12);
  assign w938[63] = |(datain[59:56] ^ 13);
  assign w938[64] = |(datain[55:52] ^ 1);
  assign w938[65] = |(datain[51:48] ^ 10);
  assign w938[66] = |(datain[47:44] ^ 8);
  assign w938[67] = |(datain[43:40] ^ 1);
  assign w938[68] = |(datain[39:36] ^ 15);
  assign w938[69] = |(datain[35:32] ^ 10);
  assign w938[70] = |(datain[31:28] ^ 1);
  assign w938[71] = |(datain[27:24] ^ 0);
  assign w938[72] = |(datain[23:20] ^ 0);
  assign w938[73] = |(datain[19:16] ^ 9);
  assign comp[938] = ~(|w938);
  wire [46-1:0] w939;
  assign w939[0] = |(datain[311:308] ^ 8);
  assign w939[1] = |(datain[307:304] ^ 14);
  assign w939[2] = |(datain[303:300] ^ 13);
  assign w939[3] = |(datain[299:296] ^ 0);
  assign w939[4] = |(datain[295:292] ^ 11);
  assign w939[5] = |(datain[291:288] ^ 12);
  assign w939[6] = |(datain[287:284] ^ 0);
  assign w939[7] = |(datain[283:280] ^ 0);
  assign w939[8] = |(datain[279:276] ^ 7);
  assign w939[9] = |(datain[275:272] ^ 12);
  assign w939[10] = |(datain[271:268] ^ 1);
  assign w939[11] = |(datain[267:264] ^ 6);
  assign w939[12] = |(datain[263:260] ^ 0);
  assign w939[13] = |(datain[259:256] ^ 7);
  assign w939[14] = |(datain[255:252] ^ 11);
  assign w939[15] = |(datain[251:248] ^ 9);
  assign w939[16] = |(datain[247:244] ^ 0);
  assign w939[17] = |(datain[243:240] ^ 15);
  assign w939[18] = |(datain[239:236] ^ 4);
  assign w939[19] = |(datain[235:232] ^ 15);
  assign w939[20] = |(datain[231:228] ^ 11);
  assign w939[21] = |(datain[227:224] ^ 3);
  assign w939[22] = |(datain[223:220] ^ 0);
  assign w939[23] = |(datain[219:216] ^ 0);
  assign w939[24] = |(datain[215:212] ^ 11);
  assign w939[25] = |(datain[211:208] ^ 10);
  assign w939[26] = |(datain[207:204] ^ 0);
  assign w939[27] = |(datain[203:200] ^ 0);
  assign w939[28] = |(datain[199:196] ^ 0);
  assign w939[29] = |(datain[195:192] ^ 1);
  assign w939[30] = |(datain[191:188] ^ 11);
  assign w939[31] = |(datain[187:184] ^ 0);
  assign w939[32] = |(datain[183:180] ^ 0);
  assign w939[33] = |(datain[179:176] ^ 3);
  assign w939[34] = |(datain[175:172] ^ 11);
  assign w939[35] = |(datain[171:168] ^ 4);
  assign w939[36] = |(datain[167:164] ^ 0);
  assign w939[37] = |(datain[163:160] ^ 2);
  assign w939[38] = |(datain[159:156] ^ 11);
  assign w939[39] = |(datain[155:152] ^ 7);
  assign w939[40] = |(datain[151:148] ^ 7);
  assign w939[41] = |(datain[147:144] ^ 12);
  assign w939[42] = |(datain[143:140] ^ 12);
  assign w939[43] = |(datain[139:136] ^ 13);
  assign w939[44] = |(datain[135:132] ^ 1);
  assign w939[45] = |(datain[131:128] ^ 3);
  assign comp[939] = ~(|w939);
  wire [76-1:0] w940;
  assign w940[0] = |(datain[311:308] ^ 11);
  assign w940[1] = |(datain[307:304] ^ 14);
  assign w940[2] = |(datain[303:300] ^ 15);
  assign w940[3] = |(datain[299:296] ^ 15);
  assign w940[4] = |(datain[295:292] ^ 7);
  assign w940[5] = |(datain[291:288] ^ 2);
  assign w940[6] = |(datain[287:284] ^ 2);
  assign w940[7] = |(datain[283:280] ^ 2);
  assign w940[8] = |(datain[279:276] ^ 8);
  assign w940[9] = |(datain[275:272] ^ 0);
  assign w940[10] = |(datain[271:268] ^ 3);
  assign w940[11] = |(datain[267:264] ^ 15);
  assign w940[12] = |(datain[263:260] ^ 15);
  assign w940[13] = |(datain[259:256] ^ 12);
  assign w940[14] = |(datain[255:252] ^ 7);
  assign w940[15] = |(datain[251:248] ^ 4);
  assign w940[16] = |(datain[247:244] ^ 1);
  assign w940[17] = |(datain[243:240] ^ 13);
  assign w940[18] = |(datain[239:236] ^ 11);
  assign w940[19] = |(datain[235:232] ^ 8);
  assign w940[20] = |(datain[231:228] ^ 0);
  assign w940[21] = |(datain[227:224] ^ 1);
  assign w940[22] = |(datain[223:220] ^ 0);
  assign w940[23] = |(datain[219:216] ^ 3);
  assign w940[24] = |(datain[215:212] ^ 11);
  assign w940[25] = |(datain[211:208] ^ 1);
  assign w940[26] = |(datain[207:204] ^ 0);
  assign w940[27] = |(datain[203:200] ^ 5);
  assign w940[28] = |(datain[199:196] ^ 5);
  assign w940[29] = |(datain[195:192] ^ 0);
  assign w940[30] = |(datain[191:188] ^ 12);
  assign w940[31] = |(datain[187:184] ^ 13);
  assign w940[32] = |(datain[183:180] ^ 1);
  assign w940[33] = |(datain[179:176] ^ 3);
  assign w940[34] = |(datain[175:172] ^ 5);
  assign w940[35] = |(datain[171:168] ^ 8);
  assign w940[36] = |(datain[167:164] ^ 8);
  assign w940[37] = |(datain[163:160] ^ 8);
  assign w940[38] = |(datain[159:156] ^ 6);
  assign w940[39] = |(datain[155:152] ^ 14);
  assign w940[40] = |(datain[151:148] ^ 0);
  assign w940[41] = |(datain[147:144] ^ 2);
  assign w940[42] = |(datain[143:140] ^ 8);
  assign w940[43] = |(datain[139:136] ^ 13);
  assign w940[44] = |(datain[135:132] ^ 11);
  assign w940[45] = |(datain[131:128] ^ 7);
  assign w940[46] = |(datain[127:124] ^ 11);
  assign w940[47] = |(datain[123:120] ^ 14);
  assign w940[48] = |(datain[119:116] ^ 0);
  assign w940[49] = |(datain[115:112] ^ 1);
  assign w940[50] = |(datain[111:108] ^ 8);
  assign w940[51] = |(datain[107:104] ^ 13);
  assign w940[52] = |(datain[103:100] ^ 11);
  assign w940[53] = |(datain[99:96] ^ 14);
  assign w940[54] = |(datain[95:92] ^ 11);
  assign w940[55] = |(datain[91:88] ^ 14);
  assign w940[56] = |(datain[87:84] ^ 0);
  assign w940[57] = |(datain[83:80] ^ 1);
  assign w940[58] = |(datain[79:76] ^ 11);
  assign w940[59] = |(datain[75:72] ^ 1);
  assign w940[60] = |(datain[71:68] ^ 2);
  assign w940[61] = |(datain[67:64] ^ 1);
  assign w940[62] = |(datain[63:60] ^ 15);
  assign w940[63] = |(datain[59:56] ^ 3);
  assign w940[64] = |(datain[55:52] ^ 10);
  assign w940[65] = |(datain[51:48] ^ 5);
  assign w940[66] = |(datain[47:44] ^ 4);
  assign w940[67] = |(datain[43:40] ^ 1);
  assign w940[68] = |(datain[39:36] ^ 8);
  assign w940[69] = |(datain[35:32] ^ 11);
  assign w940[70] = |(datain[31:28] ^ 13);
  assign w940[71] = |(datain[27:24] ^ 13);
  assign w940[72] = |(datain[23:20] ^ 12);
  assign w940[73] = |(datain[19:16] ^ 13);
  assign w940[74] = |(datain[15:12] ^ 1);
  assign w940[75] = |(datain[11:8] ^ 3);
  assign comp[940] = ~(|w940);
  wire [76-1:0] w941;
  assign w941[0] = |(datain[311:308] ^ 7);
  assign w941[1] = |(datain[307:304] ^ 12);
  assign w941[2] = |(datain[303:300] ^ 0);
  assign w941[3] = |(datain[299:296] ^ 14);
  assign w941[4] = |(datain[295:292] ^ 1);
  assign w941[5] = |(datain[291:288] ^ 15);
  assign w941[6] = |(datain[287:284] ^ 15);
  assign w941[7] = |(datain[283:280] ^ 15);
  assign w941[8] = |(datain[279:276] ^ 0);
  assign w941[9] = |(datain[275:272] ^ 14);
  assign w941[10] = |(datain[271:268] ^ 1);
  assign w941[11] = |(datain[267:264] ^ 3);
  assign w941[12] = |(datain[263:260] ^ 0);
  assign w941[13] = |(datain[259:256] ^ 4);
  assign w941[14] = |(datain[255:252] ^ 12);
  assign w941[15] = |(datain[251:248] ^ 13);
  assign w941[16] = |(datain[247:244] ^ 1);
  assign w941[17] = |(datain[243:240] ^ 2);
  assign w941[18] = |(datain[239:236] ^ 11);
  assign w941[19] = |(datain[235:232] ^ 1);
  assign w941[20] = |(datain[231:228] ^ 0);
  assign w941[21] = |(datain[227:224] ^ 10);
  assign w941[22] = |(datain[223:220] ^ 13);
  assign w941[23] = |(datain[219:216] ^ 3);
  assign w941[24] = |(datain[215:212] ^ 12);
  assign w941[25] = |(datain[211:208] ^ 8);
  assign w941[26] = |(datain[207:204] ^ 8);
  assign w941[27] = |(datain[203:200] ^ 14);
  assign w941[28] = |(datain[199:196] ^ 12);
  assign w941[29] = |(datain[195:192] ^ 0);
  assign w941[30] = |(datain[191:188] ^ 3);
  assign w941[31] = |(datain[187:184] ^ 3);
  assign w941[32] = |(datain[183:180] ^ 15);
  assign w941[33] = |(datain[179:176] ^ 15);
  assign w941[34] = |(datain[175:172] ^ 8);
  assign w941[35] = |(datain[171:168] ^ 11);
  assign w941[36] = |(datain[167:164] ^ 15);
  assign w941[37] = |(datain[163:160] ^ 4);
  assign w941[38] = |(datain[159:156] ^ 11);
  assign w941[39] = |(datain[155:152] ^ 9);
  assign w941[40] = |(datain[151:148] ^ 0);
  assign w941[41] = |(datain[147:144] ^ 0);
  assign w941[42] = |(datain[143:140] ^ 0);
  assign w941[43] = |(datain[139:136] ^ 1);
  assign w941[44] = |(datain[135:132] ^ 15);
  assign w941[45] = |(datain[131:128] ^ 3);
  assign w941[46] = |(datain[127:124] ^ 10);
  assign w941[47] = |(datain[123:120] ^ 5);
  assign w941[48] = |(datain[119:116] ^ 0);
  assign w941[49] = |(datain[115:112] ^ 6);
  assign w941[50] = |(datain[111:108] ^ 11);
  assign w941[51] = |(datain[107:104] ^ 8);
  assign w941[52] = |(datain[103:100] ^ 6);
  assign w941[53] = |(datain[99:96] ^ 3);
  assign w941[54] = |(datain[95:92] ^ 0);
  assign w941[55] = |(datain[91:88] ^ 0);
  assign w941[56] = |(datain[87:84] ^ 5);
  assign w941[57] = |(datain[83:80] ^ 0);
  assign w941[58] = |(datain[79:76] ^ 12);
  assign w941[59] = |(datain[75:72] ^ 11);
  assign w941[60] = |(datain[71:68] ^ 2);
  assign w941[61] = |(datain[67:64] ^ 14);
  assign w941[62] = |(datain[63:60] ^ 12);
  assign w941[63] = |(datain[59:56] ^ 6);
  assign w941[64] = |(datain[55:52] ^ 0);
  assign w941[65] = |(datain[51:48] ^ 6);
  assign w941[66] = |(datain[47:44] ^ 14);
  assign w941[67] = |(datain[43:40] ^ 8);
  assign w941[68] = |(datain[39:36] ^ 0);
  assign w941[69] = |(datain[35:32] ^ 1);
  assign w941[70] = |(datain[31:28] ^ 0);
  assign w941[71] = |(datain[27:24] ^ 0);
  assign w941[72] = |(datain[23:20] ^ 15);
  assign w941[73] = |(datain[19:16] ^ 15);
  assign w941[74] = |(datain[15:12] ^ 3);
  assign w941[75] = |(datain[11:8] ^ 6);
  assign comp[941] = ~(|w941);
  wire [76-1:0] w942;
  assign w942[0] = |(datain[311:308] ^ 1);
  assign w942[1] = |(datain[307:304] ^ 2);
  assign w942[2] = |(datain[303:300] ^ 2);
  assign w942[3] = |(datain[299:296] ^ 12);
  assign w942[4] = |(datain[295:292] ^ 2);
  assign w942[5] = |(datain[291:288] ^ 0);
  assign w942[6] = |(datain[287:284] ^ 13);
  assign w942[7] = |(datain[283:280] ^ 3);
  assign w942[8] = |(datain[279:276] ^ 14);
  assign w942[9] = |(datain[275:272] ^ 0);
  assign w942[10] = |(datain[271:268] ^ 11);
  assign w942[11] = |(datain[267:264] ^ 9);
  assign w942[12] = |(datain[263:260] ^ 11);
  assign w942[13] = |(datain[259:256] ^ 9);
  assign w942[14] = |(datain[255:252] ^ 0);
  assign w942[15] = |(datain[251:248] ^ 1);
  assign w942[16] = |(datain[247:244] ^ 15);
  assign w942[17] = |(datain[243:240] ^ 12);
  assign w942[18] = |(datain[239:236] ^ 8);
  assign w942[19] = |(datain[235:232] ^ 14);
  assign w942[20] = |(datain[231:228] ^ 12);
  assign w942[21] = |(datain[227:224] ^ 0);
  assign w942[22] = |(datain[223:220] ^ 15);
  assign w942[23] = |(datain[219:216] ^ 3);
  assign w942[24] = |(datain[215:212] ^ 10);
  assign w942[25] = |(datain[211:208] ^ 4);
  assign w942[26] = |(datain[207:204] ^ 11);
  assign w942[27] = |(datain[203:200] ^ 14);
  assign w942[28] = |(datain[199:196] ^ 4);
  assign w942[29] = |(datain[195:192] ^ 12);
  assign w942[30] = |(datain[191:188] ^ 0);
  assign w942[31] = |(datain[187:184] ^ 0);
  assign w942[32] = |(datain[183:180] ^ 10);
  assign w942[33] = |(datain[179:176] ^ 5);
  assign w942[34] = |(datain[175:172] ^ 10);
  assign w942[35] = |(datain[171:168] ^ 5);
  assign w942[36] = |(datain[167:164] ^ 8);
  assign w942[37] = |(datain[163:160] ^ 9);
  assign w942[38] = |(datain[159:156] ^ 4);
  assign w942[39] = |(datain[155:152] ^ 4);
  assign w942[40] = |(datain[151:148] ^ 15);
  assign w942[41] = |(datain[147:144] ^ 14);
  assign w942[42] = |(datain[143:140] ^ 12);
  assign w942[43] = |(datain[139:136] ^ 7);
  assign w942[44] = |(datain[135:132] ^ 4);
  assign w942[45] = |(datain[131:128] ^ 4);
  assign w942[46] = |(datain[127:124] ^ 15);
  assign w942[47] = |(datain[123:120] ^ 12);
  assign w942[48] = |(datain[119:116] ^ 2);
  assign w942[49] = |(datain[115:112] ^ 14);
  assign w942[50] = |(datain[111:108] ^ 7);
  assign w942[51] = |(datain[107:104] ^ 13);
  assign w942[52] = |(datain[103:100] ^ 15);
  assign w942[53] = |(datain[99:96] ^ 15);
  assign w942[54] = |(datain[95:92] ^ 0);
  assign w942[55] = |(datain[91:88] ^ 14);
  assign w942[56] = |(datain[87:84] ^ 1);
  assign w942[57] = |(datain[83:80] ^ 3);
  assign w942[58] = |(datain[79:76] ^ 0);
  assign w942[59] = |(datain[75:72] ^ 4);
  assign w942[60] = |(datain[71:68] ^ 2);
  assign w942[61] = |(datain[67:64] ^ 11);
  assign w942[62] = |(datain[63:60] ^ 12);
  assign w942[63] = |(datain[59:56] ^ 0);
  assign w942[64] = |(datain[55:52] ^ 9);
  assign w942[65] = |(datain[51:48] ^ 9);
  assign w942[66] = |(datain[47:44] ^ 12);
  assign w942[67] = |(datain[43:40] ^ 13);
  assign w942[68] = |(datain[39:36] ^ 1);
  assign w942[69] = |(datain[35:32] ^ 3);
  assign w942[70] = |(datain[31:28] ^ 12);
  assign w942[71] = |(datain[27:24] ^ 13);
  assign w942[72] = |(datain[23:20] ^ 1);
  assign w942[73] = |(datain[19:16] ^ 9);
  assign w942[74] = |(datain[15:12] ^ 9);
  assign w942[75] = |(datain[11:8] ^ 12);
  assign comp[942] = ~(|w942);
  wire [76-1:0] w943;
  assign w943[0] = |(datain[311:308] ^ 10);
  assign w943[1] = |(datain[307:304] ^ 3);
  assign w943[2] = |(datain[303:300] ^ 12);
  assign w943[3] = |(datain[299:296] ^ 4);
  assign w943[4] = |(datain[295:292] ^ 7);
  assign w943[5] = |(datain[291:288] ^ 12);
  assign w943[6] = |(datain[287:284] ^ 12);
  assign w943[7] = |(datain[283:280] ^ 1);
  assign w943[8] = |(datain[279:276] ^ 14);
  assign w943[9] = |(datain[275:272] ^ 0);
  assign w943[10] = |(datain[271:268] ^ 0);
  assign w943[11] = |(datain[267:264] ^ 6);
  assign w943[12] = |(datain[263:260] ^ 2);
  assign w943[13] = |(datain[259:256] ^ 13);
  assign w943[14] = |(datain[255:252] ^ 1);
  assign w943[15] = |(datain[251:248] ^ 10);
  assign w943[16] = |(datain[247:244] ^ 0);
  assign w943[17] = |(datain[243:240] ^ 0);
  assign w943[18] = |(datain[239:236] ^ 10);
  assign w943[19] = |(datain[235:232] ^ 3);
  assign w943[20] = |(datain[231:228] ^ 11);
  assign w943[21] = |(datain[227:224] ^ 14);
  assign w943[22] = |(datain[223:220] ^ 7);
  assign w943[23] = |(datain[219:216] ^ 12);
  assign w943[24] = |(datain[215:212] ^ 2);
  assign w943[25] = |(datain[211:208] ^ 13);
  assign w943[26] = |(datain[207:204] ^ 12);
  assign w943[27] = |(datain[203:200] ^ 3);
  assign w943[28] = |(datain[199:196] ^ 0);
  assign w943[29] = |(datain[195:192] ^ 7);
  assign w943[30] = |(datain[191:188] ^ 11);
  assign w943[31] = |(datain[187:184] ^ 9);
  assign w943[32] = |(datain[183:180] ^ 11);
  assign w943[33] = |(datain[179:176] ^ 14);
  assign w943[34] = |(datain[175:172] ^ 0);
  assign w943[35] = |(datain[171:168] ^ 1);
  assign w943[36] = |(datain[167:164] ^ 15);
  assign w943[37] = |(datain[163:160] ^ 12);
  assign w943[38] = |(datain[159:156] ^ 5);
  assign w943[39] = |(datain[155:152] ^ 0);
  assign w943[40] = |(datain[151:148] ^ 0);
  assign w943[41] = |(datain[147:144] ^ 7);
  assign w943[42] = |(datain[143:140] ^ 15);
  assign w943[43] = |(datain[139:136] ^ 3);
  assign w943[44] = |(datain[135:132] ^ 10);
  assign w943[45] = |(datain[131:128] ^ 4);
  assign w943[46] = |(datain[127:124] ^ 11);
  assign w943[47] = |(datain[123:120] ^ 14);
  assign w943[48] = |(datain[119:116] ^ 4);
  assign w943[49] = |(datain[115:112] ^ 12);
  assign w943[50] = |(datain[111:108] ^ 0);
  assign w943[51] = |(datain[107:104] ^ 0);
  assign w943[52] = |(datain[103:100] ^ 10);
  assign w943[53] = |(datain[99:96] ^ 5);
  assign w943[54] = |(datain[95:92] ^ 12);
  assign w943[55] = |(datain[91:88] ^ 7);
  assign w943[56] = |(datain[87:84] ^ 4);
  assign w943[57] = |(datain[83:80] ^ 4);
  assign w943[58] = |(datain[79:76] ^ 15);
  assign w943[59] = |(datain[75:72] ^ 14);
  assign w943[60] = |(datain[71:68] ^ 3);
  assign w943[61] = |(datain[67:64] ^ 5);
  assign w943[62] = |(datain[63:60] ^ 7);
  assign w943[63] = |(datain[59:56] ^ 13);
  assign w943[64] = |(datain[55:52] ^ 15);
  assign w943[65] = |(datain[51:48] ^ 15);
  assign w943[66] = |(datain[47:44] ^ 0);
  assign w943[67] = |(datain[43:40] ^ 14);
  assign w943[68] = |(datain[39:36] ^ 1);
  assign w943[69] = |(datain[35:32] ^ 3);
  assign w943[70] = |(datain[31:28] ^ 0);
  assign w943[71] = |(datain[27:24] ^ 4);
  assign w943[72] = |(datain[23:20] ^ 10);
  assign w943[73] = |(datain[19:16] ^ 5);
  assign w943[74] = |(datain[15:12] ^ 8);
  assign w943[75] = |(datain[11:8] ^ 9);
  assign comp[943] = ~(|w943);
  wire [74-1:0] w944;
  assign w944[0] = |(datain[311:308] ^ 3);
  assign w944[1] = |(datain[307:304] ^ 3);
  assign w944[2] = |(datain[303:300] ^ 12);
  assign w944[3] = |(datain[299:296] ^ 0);
  assign w944[4] = |(datain[295:292] ^ 15);
  assign w944[5] = |(datain[291:288] ^ 10);
  assign w944[6] = |(datain[287:284] ^ 8);
  assign w944[7] = |(datain[283:280] ^ 14);
  assign w944[8] = |(datain[279:276] ^ 13);
  assign w944[9] = |(datain[275:272] ^ 0);
  assign w944[10] = |(datain[271:268] ^ 8);
  assign w944[11] = |(datain[267:264] ^ 11);
  assign w944[12] = |(datain[263:260] ^ 14);
  assign w944[13] = |(datain[259:256] ^ 6);
  assign w944[14] = |(datain[255:252] ^ 15);
  assign w944[15] = |(datain[251:248] ^ 11);
  assign w944[16] = |(datain[247:244] ^ 8);
  assign w944[17] = |(datain[243:240] ^ 14);
  assign w944[18] = |(datain[239:236] ^ 13);
  assign w944[19] = |(datain[235:232] ^ 8);
  assign w944[20] = |(datain[231:228] ^ 8);
  assign w944[21] = |(datain[227:224] ^ 3);
  assign w944[22] = |(datain[223:220] ^ 2);
  assign w944[23] = |(datain[219:216] ^ 14);
  assign w944[24] = |(datain[215:212] ^ 1);
  assign w944[25] = |(datain[211:208] ^ 3);
  assign w944[26] = |(datain[207:204] ^ 0);
  assign w944[27] = |(datain[203:200] ^ 4);
  assign w944[28] = |(datain[199:196] ^ 0);
  assign w944[29] = |(datain[195:192] ^ 1);
  assign w944[30] = |(datain[191:188] ^ 12);
  assign w944[31] = |(datain[187:184] ^ 13);
  assign w944[32] = |(datain[183:180] ^ 1);
  assign w944[33] = |(datain[179:176] ^ 2);
  assign w944[34] = |(datain[175:172] ^ 11);
  assign w944[35] = |(datain[171:168] ^ 1);
  assign w944[36] = |(datain[167:164] ^ 0);
  assign w944[37] = |(datain[163:160] ^ 6);
  assign w944[38] = |(datain[159:156] ^ 13);
  assign w944[39] = |(datain[155:152] ^ 3);
  assign w944[40] = |(datain[151:148] ^ 14);
  assign w944[41] = |(datain[147:144] ^ 0);
  assign w944[42] = |(datain[143:140] ^ 8);
  assign w944[43] = |(datain[139:136] ^ 14);
  assign w944[44] = |(datain[135:132] ^ 12);
  assign w944[45] = |(datain[131:128] ^ 0);
  assign w944[46] = |(datain[127:124] ^ 3);
  assign w944[47] = |(datain[123:120] ^ 2);
  assign w944[48] = |(datain[119:116] ^ 15);
  assign w944[49] = |(datain[115:112] ^ 6);
  assign w944[50] = |(datain[111:108] ^ 8);
  assign w944[51] = |(datain[107:104] ^ 0);
  assign w944[52] = |(datain[103:100] ^ 15);
  assign w944[53] = |(datain[99:96] ^ 10);
  assign w944[54] = |(datain[95:92] ^ 8);
  assign w944[55] = |(datain[91:88] ^ 0);
  assign w944[56] = |(datain[87:84] ^ 7);
  assign w944[57] = |(datain[83:80] ^ 4);
  assign w944[58] = |(datain[79:76] ^ 0);
  assign w944[59] = |(datain[75:72] ^ 0);
  assign w944[60] = |(datain[71:68] ^ 3);
  assign w944[61] = |(datain[67:64] ^ 3);
  assign w944[62] = |(datain[63:60] ^ 13);
  assign w944[63] = |(datain[59:56] ^ 11);
  assign w944[64] = |(datain[55:52] ^ 11);
  assign w944[65] = |(datain[51:48] ^ 8);
  assign w944[66] = |(datain[47:44] ^ 0);
  assign w944[67] = |(datain[43:40] ^ 2);
  assign w944[68] = |(datain[39:36] ^ 0);
  assign w944[69] = |(datain[35:32] ^ 2);
  assign w944[70] = |(datain[31:28] ^ 11);
  assign w944[71] = |(datain[27:24] ^ 9);
  assign w944[72] = |(datain[23:20] ^ 0);
  assign w944[73] = |(datain[19:16] ^ 3);
  assign comp[944] = ~(|w944);
  wire [74-1:0] w945;
  assign w945[0] = |(datain[311:308] ^ 12);
  assign w945[1] = |(datain[307:304] ^ 4);
  assign w945[2] = |(datain[303:300] ^ 2);
  assign w945[3] = |(datain[299:296] ^ 14);
  assign w945[4] = |(datain[295:292] ^ 2);
  assign w945[5] = |(datain[291:288] ^ 10);
  assign w945[6] = |(datain[287:284] ^ 0);
  assign w945[7] = |(datain[283:280] ^ 0);
  assign w945[8] = |(datain[279:276] ^ 15);
  assign w945[9] = |(datain[275:272] ^ 14);
  assign w945[10] = |(datain[271:268] ^ 4);
  assign w945[11] = |(datain[267:264] ^ 6);
  assign w945[12] = |(datain[263:260] ^ 0);
  assign w945[13] = |(datain[259:256] ^ 2);
  assign w945[14] = |(datain[255:252] ^ 11);
  assign w945[15] = |(datain[251:248] ^ 4);
  assign w945[16] = |(datain[247:244] ^ 4);
  assign w945[17] = |(datain[243:240] ^ 9);
  assign w945[18] = |(datain[239:236] ^ 12);
  assign w945[19] = |(datain[235:232] ^ 13);
  assign w945[20] = |(datain[231:228] ^ 2);
  assign w945[21] = |(datain[227:224] ^ 1);
  assign w945[22] = |(datain[223:220] ^ 11);
  assign w945[23] = |(datain[219:216] ^ 15);
  assign w945[24] = |(datain[215:212] ^ 7);
  assign w945[25] = |(datain[211:208] ^ 13);
  assign w945[26] = |(datain[207:204] ^ 0);
  assign w945[27] = |(datain[203:200] ^ 3);
  assign w945[28] = |(datain[199:196] ^ 4);
  assign w945[29] = |(datain[195:192] ^ 13);
  assign w945[30] = |(datain[191:188] ^ 11);
  assign w945[31] = |(datain[187:184] ^ 4);
  assign w945[32] = |(datain[183:180] ^ 5);
  assign w945[33] = |(datain[179:176] ^ 2);
  assign w945[34] = |(datain[175:172] ^ 12);
  assign w945[35] = |(datain[171:168] ^ 13);
  assign w945[36] = |(datain[167:164] ^ 2);
  assign w945[37] = |(datain[163:160] ^ 1);
  assign w945[38] = |(datain[159:156] ^ 15);
  assign w945[39] = |(datain[155:152] ^ 12);
  assign w945[40] = |(datain[151:148] ^ 2);
  assign w945[41] = |(datain[147:144] ^ 6);
  assign w945[42] = |(datain[143:140] ^ 12);
  assign w945[43] = |(datain[139:136] ^ 5);
  assign w945[44] = |(datain[135:132] ^ 7);
  assign w945[45] = |(datain[131:128] ^ 7);
  assign w945[46] = |(datain[127:124] ^ 2);
  assign w945[47] = |(datain[123:120] ^ 2);
  assign w945[48] = |(datain[119:116] ^ 0);
  assign w945[49] = |(datain[115:112] ^ 14);
  assign w945[50] = |(datain[111:108] ^ 0);
  assign w945[51] = |(datain[107:104] ^ 7);
  assign w945[52] = |(datain[103:100] ^ 8);
  assign w945[53] = |(datain[99:96] ^ 11);
  assign w945[54] = |(datain[95:92] ^ 12);
  assign w945[55] = |(datain[91:88] ^ 7);
  assign w945[56] = |(datain[87:84] ^ 10);
  assign w945[57] = |(datain[83:80] ^ 5);
  assign w945[58] = |(datain[79:76] ^ 10);
  assign w945[59] = |(datain[75:72] ^ 5);
  assign w945[60] = |(datain[71:68] ^ 8);
  assign w945[61] = |(datain[67:64] ^ 12);
  assign w945[62] = |(datain[63:60] ^ 4);
  assign w945[63] = |(datain[59:56] ^ 12);
  assign w945[64] = |(datain[55:52] ^ 15);
  assign w945[65] = |(datain[51:48] ^ 14);
  assign w945[66] = |(datain[47:44] ^ 8);
  assign w945[67] = |(datain[43:40] ^ 9);
  assign w945[68] = |(datain[39:36] ^ 4);
  assign w945[69] = |(datain[35:32] ^ 4);
  assign w945[70] = |(datain[31:28] ^ 15);
  assign w945[71] = |(datain[27:24] ^ 12);
  assign w945[72] = |(datain[23:20] ^ 11);
  assign w945[73] = |(datain[19:16] ^ 8);
  assign comp[945] = ~(|w945);
  wire [74-1:0] w946;
  assign w946[0] = |(datain[311:308] ^ 3);
  assign w946[1] = |(datain[307:304] ^ 3);
  assign w946[2] = |(datain[303:300] ^ 12);
  assign w946[3] = |(datain[299:296] ^ 0);
  assign w946[4] = |(datain[295:292] ^ 15);
  assign w946[5] = |(datain[291:288] ^ 10);
  assign w946[6] = |(datain[287:284] ^ 11);
  assign w946[7] = |(datain[283:280] ^ 12);
  assign w946[8] = |(datain[279:276] ^ 0);
  assign w946[9] = |(datain[275:272] ^ 0);
  assign w946[10] = |(datain[271:268] ^ 7);
  assign w946[11] = |(datain[267:264] ^ 12);
  assign w946[12] = |(datain[263:260] ^ 8);
  assign w946[13] = |(datain[259:256] ^ 14);
  assign w946[14] = |(datain[255:252] ^ 13);
  assign w946[15] = |(datain[251:248] ^ 0);
  assign w946[16] = |(datain[247:244] ^ 15);
  assign w946[17] = |(datain[243:240] ^ 11);
  assign w946[18] = |(datain[239:236] ^ 3);
  assign w946[19] = |(datain[235:232] ^ 3);
  assign w946[20] = |(datain[231:228] ^ 15);
  assign w946[21] = |(datain[227:224] ^ 15);
  assign w946[22] = |(datain[223:220] ^ 11);
  assign w946[23] = |(datain[219:216] ^ 14);
  assign w946[24] = |(datain[215:212] ^ 5);
  assign w946[25] = |(datain[211:208] ^ 0);
  assign w946[26] = |(datain[207:204] ^ 6);
  assign w946[27] = |(datain[203:200] ^ 1);
  assign w946[28] = |(datain[199:196] ^ 8);
  assign w946[29] = |(datain[195:192] ^ 14);
  assign w946[30] = |(datain[191:188] ^ 13);
  assign w946[31] = |(datain[187:184] ^ 8);
  assign w946[32] = |(datain[183:180] ^ 8);
  assign w946[33] = |(datain[179:176] ^ 1);
  assign w946[34] = |(datain[175:172] ^ 15);
  assign w946[35] = |(datain[171:168] ^ 6);
  assign w946[36] = |(datain[167:164] ^ 4);
  assign w946[37] = |(datain[163:160] ^ 3);
  assign w946[38] = |(datain[159:156] ^ 6);
  assign w946[39] = |(datain[155:152] ^ 5);
  assign w946[40] = |(datain[151:148] ^ 8);
  assign w946[41] = |(datain[147:144] ^ 3);
  assign w946[42] = |(datain[143:140] ^ 2);
  assign w946[43] = |(datain[139:136] ^ 12);
  assign w946[44] = |(datain[135:132] ^ 0);
  assign w946[45] = |(datain[131:128] ^ 4);
  assign w946[46] = |(datain[127:124] ^ 8);
  assign w946[47] = |(datain[123:120] ^ 11);
  assign w946[48] = |(datain[119:116] ^ 0);
  assign w946[49] = |(datain[115:112] ^ 4);
  assign w946[50] = |(datain[111:108] ^ 12);
  assign w946[51] = |(datain[107:104] ^ 1);
  assign w946[52] = |(datain[103:100] ^ 14);
  assign w946[53] = |(datain[99:96] ^ 0);
  assign w946[54] = |(datain[95:92] ^ 0);
  assign w946[55] = |(datain[91:88] ^ 6);
  assign w946[56] = |(datain[87:84] ^ 11);
  assign w946[57] = |(datain[83:80] ^ 14);
  assign w946[58] = |(datain[79:76] ^ 0);
  assign w946[59] = |(datain[75:72] ^ 0);
  assign w946[60] = |(datain[71:68] ^ 7);
  assign w946[61] = |(datain[67:64] ^ 12);
  assign w946[62] = |(datain[63:60] ^ 8);
  assign w946[63] = |(datain[59:56] ^ 14);
  assign w946[64] = |(datain[55:52] ^ 12);
  assign w946[65] = |(datain[51:48] ^ 0);
  assign w946[66] = |(datain[47:44] ^ 0);
  assign w946[67] = |(datain[43:40] ^ 14);
  assign w946[68] = |(datain[39:36] ^ 1);
  assign w946[69] = |(datain[35:32] ^ 15);
  assign w946[70] = |(datain[31:28] ^ 15);
  assign w946[71] = |(datain[27:24] ^ 3);
  assign w946[72] = |(datain[23:20] ^ 10);
  assign w946[73] = |(datain[19:16] ^ 4);
  assign comp[946] = ~(|w946);
  wire [76-1:0] w947;
  assign w947[0] = |(datain[311:308] ^ 15);
  assign w947[1] = |(datain[307:304] ^ 8);
  assign w947[2] = |(datain[303:300] ^ 12);
  assign w947[3] = |(datain[299:296] ^ 3);
  assign w947[4] = |(datain[295:292] ^ 15);
  assign w947[5] = |(datain[291:288] ^ 9);
  assign w947[6] = |(datain[287:284] ^ 12);
  assign w947[7] = |(datain[283:280] ^ 3);
  assign w947[8] = |(datain[279:276] ^ 5);
  assign w947[9] = |(datain[275:272] ^ 0);
  assign w947[10] = |(datain[271:268] ^ 5);
  assign w947[11] = |(datain[267:264] ^ 3);
  assign w947[12] = |(datain[263:260] ^ 5);
  assign w947[13] = |(datain[259:256] ^ 1);
  assign w947[14] = |(datain[255:252] ^ 5);
  assign w947[15] = |(datain[251:248] ^ 2);
  assign w947[16] = |(datain[247:244] ^ 3);
  assign w947[17] = |(datain[243:240] ^ 10);
  assign w947[18] = |(datain[239:236] ^ 1);
  assign w947[19] = |(datain[235:232] ^ 6);
  assign w947[20] = |(datain[231:228] ^ 7);
  assign w947[21] = |(datain[227:224] ^ 7);
  assign w947[22] = |(datain[223:220] ^ 0);
  assign w947[23] = |(datain[219:216] ^ 1);
  assign w947[24] = |(datain[215:212] ^ 8);
  assign w947[25] = |(datain[211:208] ^ 8);
  assign w947[26] = |(datain[207:204] ^ 1);
  assign w947[27] = |(datain[203:200] ^ 6);
  assign w947[28] = |(datain[199:196] ^ 7);
  assign w947[29] = |(datain[195:192] ^ 7);
  assign w947[30] = |(datain[191:188] ^ 0);
  assign w947[31] = |(datain[187:184] ^ 1);
  assign w947[32] = |(datain[183:180] ^ 7);
  assign w947[33] = |(datain[179:176] ^ 5);
  assign w947[34] = |(datain[175:172] ^ 1);
  assign w947[35] = |(datain[171:168] ^ 3);
  assign w947[36] = |(datain[167:164] ^ 3);
  assign w947[37] = |(datain[163:160] ^ 3);
  assign w947[38] = |(datain[159:156] ^ 12);
  assign w947[39] = |(datain[155:152] ^ 0);
  assign w947[40] = |(datain[151:148] ^ 12);
  assign w947[41] = |(datain[147:144] ^ 13);
  assign w947[42] = |(datain[143:140] ^ 1);
  assign w947[43] = |(datain[139:136] ^ 10);
  assign w947[44] = |(datain[135:132] ^ 8);
  assign w947[45] = |(datain[131:128] ^ 11);
  assign w947[46] = |(datain[127:124] ^ 12);
  assign w947[47] = |(datain[123:120] ^ 2);
  assign w947[48] = |(datain[119:116] ^ 2);
  assign w947[49] = |(datain[115:112] ^ 11);
  assign w947[50] = |(datain[111:108] ^ 0);
  assign w947[51] = |(datain[107:104] ^ 6);
  assign w947[52] = |(datain[103:100] ^ 7);
  assign w947[53] = |(datain[99:96] ^ 5);
  assign w947[54] = |(datain[95:92] ^ 0);
  assign w947[55] = |(datain[91:88] ^ 1);
  assign w947[56] = |(datain[87:84] ^ 8);
  assign w947[57] = |(datain[83:80] ^ 9);
  assign w947[58] = |(datain[79:76] ^ 1);
  assign w947[59] = |(datain[75:72] ^ 6);
  assign w947[60] = |(datain[71:68] ^ 7);
  assign w947[61] = |(datain[67:64] ^ 5);
  assign w947[62] = |(datain[63:60] ^ 0);
  assign w947[63] = |(datain[59:56] ^ 1);
  assign w947[64] = |(datain[55:52] ^ 3);
  assign w947[65] = |(datain[51:48] ^ 13);
  assign w947[66] = |(datain[47:44] ^ 3);
  assign w947[67] = |(datain[43:40] ^ 6);
  assign w947[68] = |(datain[39:36] ^ 0);
  assign w947[69] = |(datain[35:32] ^ 0);
  assign w947[70] = |(datain[31:28] ^ 7);
  assign w947[71] = |(datain[27:24] ^ 2);
  assign w947[72] = |(datain[23:20] ^ 0);
  assign w947[73] = |(datain[19:16] ^ 7);
  assign w947[74] = |(datain[15:12] ^ 5);
  assign w947[75] = |(datain[11:8] ^ 10);
  assign comp[947] = ~(|w947);
  wire [74-1:0] w948;
  assign w948[0] = |(datain[311:308] ^ 13);
  assign w948[1] = |(datain[307:304] ^ 8);
  assign w948[2] = |(datain[303:300] ^ 0);
  assign w948[3] = |(datain[299:296] ^ 5);
  assign w948[4] = |(datain[295:292] ^ 14);
  assign w948[5] = |(datain[291:288] ^ 10);
  assign w948[6] = |(datain[287:284] ^ 7);
  assign w948[7] = |(datain[283:280] ^ 4);
  assign w948[8] = |(datain[279:276] ^ 4);
  assign w948[9] = |(datain[275:272] ^ 1);
  assign w948[10] = |(datain[271:268] ^ 6);
  assign w948[11] = |(datain[267:264] ^ 0);
  assign w948[12] = |(datain[263:260] ^ 11);
  assign w948[13] = |(datain[259:256] ^ 14);
  assign w948[14] = |(datain[255:252] ^ 0);
  assign w948[15] = |(datain[251:248] ^ 5);
  assign w948[16] = |(datain[247:244] ^ 0);
  assign w948[17] = |(datain[243:240] ^ 0);
  assign w948[18] = |(datain[239:236] ^ 11);
  assign w948[19] = |(datain[235:232] ^ 9);
  assign w948[20] = |(datain[231:228] ^ 1);
  assign w948[21] = |(datain[227:224] ^ 11);
  assign w948[22] = |(datain[223:220] ^ 0);
  assign w948[23] = |(datain[219:216] ^ 0);
  assign w948[24] = |(datain[215:212] ^ 2);
  assign w948[25] = |(datain[211:208] ^ 6);
  assign w948[26] = |(datain[207:204] ^ 8);
  assign w948[27] = |(datain[203:200] ^ 10);
  assign w948[28] = |(datain[199:196] ^ 4);
  assign w948[29] = |(datain[195:192] ^ 7);
  assign w948[30] = |(datain[191:188] ^ 0);
  assign w948[31] = |(datain[187:184] ^ 5);
  assign w948[32] = |(datain[183:180] ^ 2);
  assign w948[33] = |(datain[179:176] ^ 14);
  assign w948[34] = |(datain[175:172] ^ 8);
  assign w948[35] = |(datain[171:168] ^ 8);
  assign w948[36] = |(datain[167:164] ^ 0);
  assign w948[37] = |(datain[163:160] ^ 4);
  assign w948[38] = |(datain[159:156] ^ 4);
  assign w948[39] = |(datain[155:152] ^ 6);
  assign w948[40] = |(datain[151:148] ^ 4);
  assign w948[41] = |(datain[147:144] ^ 3);
  assign w948[42] = |(datain[143:140] ^ 14);
  assign w948[43] = |(datain[139:136] ^ 2);
  assign w948[44] = |(datain[135:132] ^ 15);
  assign w948[45] = |(datain[131:128] ^ 5);
  assign w948[46] = |(datain[127:124] ^ 2);
  assign w948[47] = |(datain[123:120] ^ 14);
  assign w948[48] = |(datain[119:116] ^ 8);
  assign w948[49] = |(datain[115:112] ^ 8);
  assign w948[50] = |(datain[111:108] ^ 0);
  assign w948[51] = |(datain[107:104] ^ 14);
  assign w948[52] = |(datain[103:100] ^ 0);
  assign w948[53] = |(datain[99:96] ^ 4);
  assign w948[54] = |(datain[95:92] ^ 0);
  assign w948[55] = |(datain[91:88] ^ 0);
  assign w948[56] = |(datain[87:84] ^ 0);
  assign w948[57] = |(datain[83:80] ^ 6);
  assign w948[58] = |(datain[79:76] ^ 0);
  assign w948[59] = |(datain[75:72] ^ 14);
  assign w948[60] = |(datain[71:68] ^ 0);
  assign w948[61] = |(datain[67:64] ^ 7);
  assign w948[62] = |(datain[63:60] ^ 2);
  assign w948[63] = |(datain[59:56] ^ 14);
  assign w948[64] = |(datain[55:52] ^ 8);
  assign w948[65] = |(datain[51:48] ^ 11);
  assign w948[66] = |(datain[47:44] ^ 2);
  assign w948[67] = |(datain[43:40] ^ 14);
  assign w948[68] = |(datain[39:36] ^ 0);
  assign w948[69] = |(datain[35:32] ^ 3);
  assign w948[70] = |(datain[31:28] ^ 0);
  assign w948[71] = |(datain[27:24] ^ 0);
  assign w948[72] = |(datain[23:20] ^ 2);
  assign w948[73] = |(datain[19:16] ^ 14);
  assign comp[948] = ~(|w948);
  wire [76-1:0] w949;
  assign w949[0] = |(datain[311:308] ^ 7);
  assign w949[1] = |(datain[307:304] ^ 12);
  assign w949[2] = |(datain[303:300] ^ 11);
  assign w949[3] = |(datain[299:296] ^ 11);
  assign w949[4] = |(datain[295:292] ^ 0);
  assign w949[5] = |(datain[291:288] ^ 2);
  assign w949[6] = |(datain[287:284] ^ 0);
  assign w949[7] = |(datain[283:280] ^ 3);
  assign w949[8] = |(datain[279:276] ^ 3);
  assign w949[9] = |(datain[275:272] ^ 3);
  assign w949[10] = |(datain[271:268] ^ 12);
  assign w949[11] = |(datain[267:264] ^ 0);
  assign w949[12] = |(datain[263:260] ^ 8);
  assign w949[13] = |(datain[259:256] ^ 14);
  assign w949[14] = |(datain[255:252] ^ 12);
  assign w949[15] = |(datain[251:248] ^ 0);
  assign w949[16] = |(datain[247:244] ^ 15);
  assign w949[17] = |(datain[243:240] ^ 10);
  assign w949[18] = |(datain[239:236] ^ 8);
  assign w949[19] = |(datain[235:232] ^ 14);
  assign w949[20] = |(datain[231:228] ^ 13);
  assign w949[21] = |(datain[227:224] ^ 0);
  assign w949[22] = |(datain[223:220] ^ 8);
  assign w949[23] = |(datain[219:216] ^ 11);
  assign w949[24] = |(datain[215:212] ^ 14);
  assign w949[25] = |(datain[211:208] ^ 6);
  assign w949[26] = |(datain[207:204] ^ 15);
  assign w949[27] = |(datain[203:200] ^ 11);
  assign w949[28] = |(datain[199:196] ^ 8);
  assign w949[29] = |(datain[195:192] ^ 14);
  assign w949[30] = |(datain[191:188] ^ 13);
  assign w949[31] = |(datain[187:184] ^ 8);
  assign w949[32] = |(datain[183:180] ^ 15);
  assign w949[33] = |(datain[179:176] ^ 15);
  assign w949[34] = |(datain[175:172] ^ 8);
  assign w949[35] = |(datain[171:168] ^ 15);
  assign w949[36] = |(datain[167:164] ^ 1);
  assign w949[37] = |(datain[163:160] ^ 1);
  assign w949[38] = |(datain[159:156] ^ 0);
  assign w949[39] = |(datain[155:152] ^ 1);
  assign w949[40] = |(datain[151:148] ^ 8);
  assign w949[41] = |(datain[147:144] ^ 11);
  assign w949[42] = |(datain[143:140] ^ 8);
  assign w949[43] = |(datain[139:136] ^ 7);
  assign w949[44] = |(datain[135:132] ^ 1);
  assign w949[45] = |(datain[131:128] ^ 1);
  assign w949[46] = |(datain[127:124] ^ 0);
  assign w949[47] = |(datain[123:120] ^ 1);
  assign w949[48] = |(datain[119:116] ^ 12);
  assign w949[49] = |(datain[115:112] ^ 1);
  assign w949[50] = |(datain[111:108] ^ 14);
  assign w949[51] = |(datain[107:104] ^ 0);
  assign w949[52] = |(datain[103:100] ^ 0);
  assign w949[53] = |(datain[99:96] ^ 6);
  assign w949[54] = |(datain[95:92] ^ 8);
  assign w949[55] = |(datain[91:88] ^ 14);
  assign w949[56] = |(datain[87:84] ^ 12);
  assign w949[57] = |(datain[83:80] ^ 0);
  assign w949[58] = |(datain[79:76] ^ 11);
  assign w949[59] = |(datain[75:72] ^ 8);
  assign w949[60] = |(datain[71:68] ^ 0);
  assign w949[61] = |(datain[67:64] ^ 0);
  assign w949[62] = |(datain[63:60] ^ 0);
  assign w949[63] = |(datain[59:56] ^ 2);
  assign w949[64] = |(datain[55:52] ^ 9);
  assign w949[65] = |(datain[51:48] ^ 1);
  assign w949[66] = |(datain[47:44] ^ 8);
  assign w949[67] = |(datain[43:40] ^ 0);
  assign w949[68] = |(datain[39:36] ^ 15);
  assign w949[69] = |(datain[35:32] ^ 10);
  assign w949[70] = |(datain[31:28] ^ 8);
  assign w949[71] = |(datain[27:24] ^ 0);
  assign w949[72] = |(datain[23:20] ^ 7);
  assign w949[73] = |(datain[19:16] ^ 4);
  assign w949[74] = |(datain[15:12] ^ 0);
  assign w949[75] = |(datain[11:8] ^ 3);
  assign comp[949] = ~(|w949);
  wire [76-1:0] w950;
  assign w950[0] = |(datain[311:308] ^ 10);
  assign w950[1] = |(datain[307:304] ^ 1);
  assign w950[2] = |(datain[303:300] ^ 1);
  assign w950[3] = |(datain[299:296] ^ 3);
  assign w950[4] = |(datain[295:292] ^ 0);
  assign w950[5] = |(datain[291:288] ^ 4);
  assign w950[6] = |(datain[287:284] ^ 13);
  assign w950[7] = |(datain[283:280] ^ 3);
  assign w950[8] = |(datain[279:276] ^ 14);
  assign w950[9] = |(datain[275:272] ^ 0);
  assign w950[10] = |(datain[271:268] ^ 2);
  assign w950[11] = |(datain[267:264] ^ 13);
  assign w950[12] = |(datain[263:260] ^ 14);
  assign w950[13] = |(datain[259:256] ^ 0);
  assign w950[14] = |(datain[255:252] ^ 0);
  assign w950[15] = |(datain[251:248] ^ 7);
  assign w950[16] = |(datain[247:244] ^ 8);
  assign w950[17] = |(datain[243:240] ^ 14);
  assign w950[18] = |(datain[239:236] ^ 12);
  assign w950[19] = |(datain[235:232] ^ 0);
  assign w950[20] = |(datain[231:228] ^ 8);
  assign w950[21] = |(datain[227:224] ^ 3);
  assign w950[22] = |(datain[223:220] ^ 2);
  assign w950[23] = |(datain[219:216] ^ 14);
  assign w950[24] = |(datain[215:212] ^ 1);
  assign w950[25] = |(datain[211:208] ^ 3);
  assign w950[26] = |(datain[207:204] ^ 0);
  assign w950[27] = |(datain[203:200] ^ 4);
  assign w950[28] = |(datain[199:196] ^ 0);
  assign w950[29] = |(datain[195:192] ^ 3);
  assign w950[30] = |(datain[191:188] ^ 11);
  assign w950[31] = |(datain[187:184] ^ 14);
  assign w950[32] = |(datain[183:180] ^ 0);
  assign w950[33] = |(datain[179:176] ^ 0);
  assign w950[34] = |(datain[175:172] ^ 7);
  assign w950[35] = |(datain[171:168] ^ 12);
  assign w950[36] = |(datain[167:164] ^ 8);
  assign w950[37] = |(datain[163:160] ^ 11);
  assign w950[38] = |(datain[159:156] ^ 15);
  assign w950[39] = |(datain[155:152] ^ 14);
  assign w950[40] = |(datain[151:148] ^ 11);
  assign w950[41] = |(datain[147:144] ^ 9);
  assign w950[42] = |(datain[143:140] ^ 0);
  assign w950[43] = |(datain[139:136] ^ 0);
  assign w950[44] = |(datain[135:132] ^ 0);
  assign w950[45] = |(datain[131:128] ^ 1);
  assign w950[46] = |(datain[127:124] ^ 15);
  assign w950[47] = |(datain[123:120] ^ 3);
  assign w950[48] = |(datain[119:116] ^ 10);
  assign w950[49] = |(datain[115:112] ^ 5);
  assign w950[50] = |(datain[111:108] ^ 0);
  assign w950[51] = |(datain[107:104] ^ 6);
  assign w950[52] = |(datain[103:100] ^ 11);
  assign w950[53] = |(datain[99:96] ^ 8);
  assign w950[54] = |(datain[95:92] ^ 7);
  assign w950[55] = |(datain[91:88] ^ 0);
  assign w950[56] = |(datain[87:84] ^ 7);
  assign w950[57] = |(datain[83:80] ^ 12);
  assign w950[58] = |(datain[79:76] ^ 5);
  assign w950[59] = |(datain[75:72] ^ 0);
  assign w950[60] = |(datain[71:68] ^ 12);
  assign w950[61] = |(datain[67:64] ^ 11);
  assign w950[62] = |(datain[63:60] ^ 0);
  assign w950[63] = |(datain[59:56] ^ 6);
  assign w950[64] = |(datain[55:52] ^ 1);
  assign w950[65] = |(datain[51:48] ^ 15);
  assign w950[66] = |(datain[47:44] ^ 11);
  assign w950[67] = |(datain[43:40] ^ 11);
  assign w950[68] = |(datain[39:36] ^ 0);
  assign w950[69] = |(datain[35:32] ^ 0);
  assign w950[70] = |(datain[31:28] ^ 7);
  assign w950[71] = |(datain[27:24] ^ 2);
  assign w950[72] = |(datain[23:20] ^ 8);
  assign w950[73] = |(datain[19:16] ^ 11);
  assign w950[74] = |(datain[15:12] ^ 0);
  assign w950[75] = |(datain[11:8] ^ 14);
  assign comp[950] = ~(|w950);
  wire [74-1:0] w951;
  assign w951[0] = |(datain[311:308] ^ 3);
  assign w951[1] = |(datain[307:304] ^ 11);
  assign w951[2] = |(datain[303:300] ^ 0);
  assign w951[3] = |(datain[299:296] ^ 6);
  assign w951[4] = |(datain[295:292] ^ 2);
  assign w951[5] = |(datain[291:288] ^ 3);
  assign w951[6] = |(datain[287:284] ^ 0);
  assign w951[7] = |(datain[283:280] ^ 3);
  assign w951[8] = |(datain[279:276] ^ 7);
  assign w951[9] = |(datain[275:272] ^ 4);
  assign w951[10] = |(datain[271:268] ^ 2);
  assign w951[11] = |(datain[267:264] ^ 13);
  assign w951[12] = |(datain[263:260] ^ 14);
  assign w951[13] = |(datain[259:256] ^ 8);
  assign w951[14] = |(datain[255:252] ^ 5);
  assign w951[15] = |(datain[251:248] ^ 13);
  assign w951[16] = |(datain[247:244] ^ 0);
  assign w951[17] = |(datain[243:240] ^ 0);
  assign w951[18] = |(datain[239:236] ^ 12);
  assign w951[19] = |(datain[235:232] ^ 6);
  assign w951[20] = |(datain[231:228] ^ 0);
  assign w951[21] = |(datain[227:224] ^ 6);
  assign w951[22] = |(datain[223:220] ^ 11);
  assign w951[23] = |(datain[219:216] ^ 15);
  assign w951[24] = |(datain[215:212] ^ 0);
  assign w951[25] = |(datain[211:208] ^ 0);
  assign w951[26] = |(datain[207:204] ^ 0);
  assign w951[27] = |(datain[203:200] ^ 0);
  assign w951[28] = |(datain[199:196] ^ 8);
  assign w951[29] = |(datain[195:192] ^ 0);
  assign w951[30] = |(datain[191:188] ^ 15);
  assign w951[31] = |(datain[187:184] ^ 10);
  assign w951[32] = |(datain[183:180] ^ 8);
  assign w951[33] = |(datain[179:176] ^ 0);
  assign w951[34] = |(datain[175:172] ^ 7);
  assign w951[35] = |(datain[171:168] ^ 4);
  assign w951[36] = |(datain[167:164] ^ 1);
  assign w951[37] = |(datain[163:160] ^ 9);
  assign w951[38] = |(datain[159:156] ^ 11);
  assign w951[39] = |(datain[155:152] ^ 4);
  assign w951[40] = |(datain[151:148] ^ 0);
  assign w951[41] = |(datain[147:144] ^ 3);
  assign w951[42] = |(datain[143:140] ^ 11);
  assign w951[43] = |(datain[139:136] ^ 11);
  assign w951[44] = |(datain[135:132] ^ 0);
  assign w951[45] = |(datain[131:128] ^ 0);
  assign w951[46] = |(datain[127:124] ^ 0);
  assign w951[47] = |(datain[123:120] ^ 2);
  assign w951[48] = |(datain[119:116] ^ 11);
  assign w951[49] = |(datain[115:112] ^ 1);
  assign w951[50] = |(datain[111:108] ^ 0);
  assign w951[51] = |(datain[107:104] ^ 3);
  assign w951[52] = |(datain[103:100] ^ 11);
  assign w951[53] = |(datain[99:96] ^ 6);
  assign w951[54] = |(datain[95:92] ^ 0);
  assign w951[55] = |(datain[91:88] ^ 1);
  assign w951[56] = |(datain[87:84] ^ 8);
  assign w951[57] = |(datain[83:80] ^ 0);
  assign w951[58] = |(datain[79:76] ^ 3);
  assign w951[59] = |(datain[75:72] ^ 14);
  assign w951[60] = |(datain[71:68] ^ 1);
  assign w951[61] = |(datain[67:64] ^ 5);
  assign w951[62] = |(datain[63:60] ^ 0);
  assign w951[63] = |(datain[59:56] ^ 2);
  assign w951[64] = |(datain[55:52] ^ 15);
  assign w951[65] = |(datain[51:48] ^ 13);
  assign w951[66] = |(datain[47:44] ^ 7);
  assign w951[67] = |(datain[43:40] ^ 4);
  assign w951[68] = |(datain[39:36] ^ 0);
  assign w951[69] = |(datain[35:32] ^ 2);
  assign w951[70] = |(datain[31:28] ^ 11);
  assign w951[71] = |(datain[27:24] ^ 1);
  assign w951[72] = |(datain[23:20] ^ 0);
  assign w951[73] = |(datain[19:16] ^ 14);
  assign comp[951] = ~(|w951);
  wire [42-1:0] w952;
  assign w952[0] = |(datain[311:308] ^ 13);
  assign w952[1] = |(datain[307:304] ^ 8);
  assign w952[2] = |(datain[303:300] ^ 10);
  assign w952[3] = |(datain[299:296] ^ 1);
  assign w952[4] = |(datain[295:292] ^ 6);
  assign w952[5] = |(datain[291:288] ^ 13);
  assign w952[6] = |(datain[287:284] ^ 0);
  assign w952[7] = |(datain[283:280] ^ 4);
  assign w952[8] = |(datain[279:276] ^ 2);
  assign w952[9] = |(datain[275:272] ^ 5);
  assign w952[10] = |(datain[271:268] ^ 8);
  assign w952[11] = |(datain[267:264] ^ 15);
  assign w952[12] = |(datain[263:260] ^ 1);
  assign w952[13] = |(datain[259:256] ^ 7);
  assign w952[14] = |(datain[255:252] ^ 7);
  assign w952[15] = |(datain[251:248] ^ 5);
  assign w952[16] = |(datain[247:244] ^ 1);
  assign w952[17] = |(datain[243:240] ^ 0);
  assign w952[18] = |(datain[239:236] ^ 14);
  assign w952[19] = |(datain[235:232] ^ 8);
  assign w952[20] = |(datain[231:228] ^ 11);
  assign w952[21] = |(datain[227:224] ^ 8);
  assign w952[22] = |(datain[223:220] ^ 0);
  assign w952[23] = |(datain[219:216] ^ 0);
  assign w952[24] = |(datain[215:212] ^ 5);
  assign w952[25] = |(datain[211:208] ^ 0);
  assign w952[26] = |(datain[207:204] ^ 14);
  assign w952[27] = |(datain[203:200] ^ 8);
  assign w952[28] = |(datain[199:196] ^ 9);
  assign w952[29] = |(datain[195:192] ^ 15);
  assign w952[30] = |(datain[191:188] ^ 0);
  assign w952[31] = |(datain[187:184] ^ 0);
  assign w952[32] = |(datain[183:180] ^ 8);
  assign w952[33] = |(datain[179:176] ^ 1);
  assign w952[34] = |(datain[175:172] ^ 15);
  assign w952[35] = |(datain[171:168] ^ 1);
  assign w952[36] = |(datain[167:164] ^ 12);
  assign w952[37] = |(datain[163:160] ^ 0);
  assign w952[38] = |(datain[159:156] ^ 15);
  assign w952[39] = |(datain[155:152] ^ 15);
  assign w952[40] = |(datain[151:148] ^ 13);
  assign w952[41] = |(datain[147:144] ^ 1);
  assign comp[952] = ~(|w952);
  wire [60-1:0] w953;
  assign w953[0] = |(datain[311:308] ^ 15);
  assign w953[1] = |(datain[307:304] ^ 6);
  assign w953[2] = |(datain[303:300] ^ 4);
  assign w953[3] = |(datain[299:296] ^ 8);
  assign w953[4] = |(datain[295:292] ^ 5);
  assign w953[5] = |(datain[291:288] ^ 10);
  assign w953[6] = |(datain[287:284] ^ 8);
  assign w953[7] = |(datain[283:280] ^ 8);
  assign w953[8] = |(datain[279:276] ^ 12);
  assign w953[9] = |(datain[275:272] ^ 5);
  assign w953[10] = |(datain[271:268] ^ 11);
  assign w953[11] = |(datain[267:264] ^ 1);
  assign w953[12] = |(datain[263:260] ^ 0);
  assign w953[13] = |(datain[259:256] ^ 1);
  assign w953[14] = |(datain[255:252] ^ 3);
  assign w953[15] = |(datain[251:248] ^ 3);
  assign w953[16] = |(datain[247:244] ^ 13);
  assign w953[17] = |(datain[243:240] ^ 11);
  assign w953[18] = |(datain[239:236] ^ 11);
  assign w953[19] = |(datain[235:232] ^ 8);
  assign w953[20] = |(datain[231:228] ^ 0);
  assign w953[21] = |(datain[227:224] ^ 3);
  assign w953[22] = |(datain[223:220] ^ 0);
  assign w953[23] = |(datain[219:216] ^ 2);
  assign w953[24] = |(datain[215:212] ^ 11);
  assign w953[25] = |(datain[211:208] ^ 6);
  assign w953[26] = |(datain[207:204] ^ 0);
  assign w953[27] = |(datain[203:200] ^ 1);
  assign w953[28] = |(datain[199:196] ^ 8);
  assign w953[29] = |(datain[195:192] ^ 10);
  assign w953[30] = |(datain[191:188] ^ 1);
  assign w953[31] = |(datain[187:184] ^ 6);
  assign w953[32] = |(datain[183:180] ^ 9);
  assign w953[33] = |(datain[179:176] ^ 0);
  assign w953[34] = |(datain[175:172] ^ 7);
  assign w953[35] = |(datain[171:168] ^ 12);
  assign w953[36] = |(datain[167:164] ^ 12);
  assign w953[37] = |(datain[163:160] ^ 13);
  assign w953[38] = |(datain[159:156] ^ 1);
  assign w953[39] = |(datain[155:152] ^ 3);
  assign w953[40] = |(datain[151:148] ^ 8);
  assign w953[41] = |(datain[147:144] ^ 12);
  assign w953[42] = |(datain[143:140] ^ 12);
  assign w953[43] = |(datain[139:136] ^ 0);
  assign w953[44] = |(datain[135:132] ^ 0);
  assign w953[45] = |(datain[131:128] ^ 5);
  assign w953[46] = |(datain[127:124] ^ 2);
  assign w953[47] = |(datain[123:120] ^ 0);
  assign w953[48] = |(datain[119:116] ^ 0);
  assign w953[49] = |(datain[115:112] ^ 0);
  assign w953[50] = |(datain[111:108] ^ 5);
  assign w953[51] = |(datain[107:104] ^ 0);
  assign w953[52] = |(datain[103:100] ^ 6);
  assign w953[53] = |(datain[99:96] ^ 8);
  assign w953[54] = |(datain[95:92] ^ 0);
  assign w953[55] = |(datain[91:88] ^ 5);
  assign w953[56] = |(datain[87:84] ^ 0);
  assign w953[57] = |(datain[83:80] ^ 3);
  assign w953[58] = |(datain[79:76] ^ 12);
  assign w953[59] = |(datain[75:72] ^ 11);
  assign comp[953] = ~(|w953);
  wire [70-1:0] w954;
  assign w954[0] = |(datain[311:308] ^ 8);
  assign w954[1] = |(datain[307:304] ^ 11);
  assign w954[2] = |(datain[303:300] ^ 14);
  assign w954[3] = |(datain[299:296] ^ 12);
  assign w954[4] = |(datain[295:292] ^ 12);
  assign w954[5] = |(datain[291:288] ^ 7);
  assign w954[6] = |(datain[287:284] ^ 4);
  assign w954[7] = |(datain[283:280] ^ 6);
  assign w954[8] = |(datain[279:276] ^ 0);
  assign w954[9] = |(datain[275:272] ^ 2);
  assign w954[10] = |(datain[271:268] ^ 0);
  assign w954[11] = |(datain[267:264] ^ 0);
  assign w954[12] = |(datain[263:260] ^ 0);
  assign w954[13] = |(datain[259:256] ^ 0);
  assign w954[14] = |(datain[255:252] ^ 5);
  assign w954[15] = |(datain[251:248] ^ 13);
  assign w954[16] = |(datain[247:244] ^ 1);
  assign w954[17] = |(datain[243:240] ^ 15);
  assign w954[18] = |(datain[239:236] ^ 10);
  assign w954[19] = |(datain[235:232] ^ 0);
  assign w954[20] = |(datain[231:228] ^ 3);
  assign w954[21] = |(datain[227:224] ^ 15);
  assign w954[22] = |(datain[223:220] ^ 0);
  assign w954[23] = |(datain[219:216] ^ 4);
  assign w954[24] = |(datain[215:212] ^ 5);
  assign w954[25] = |(datain[211:208] ^ 1);
  assign w954[26] = |(datain[207:204] ^ 11);
  assign w954[27] = |(datain[203:200] ^ 1);
  assign w954[28] = |(datain[199:196] ^ 0);
  assign w954[29] = |(datain[195:192] ^ 4);
  assign w954[30] = |(datain[191:188] ^ 13);
  assign w954[31] = |(datain[187:184] ^ 2);
  assign w954[32] = |(datain[183:180] ^ 14);
  assign w954[33] = |(datain[179:176] ^ 0);
  assign w954[34] = |(datain[175:172] ^ 5);
  assign w954[35] = |(datain[171:168] ^ 9);
  assign w954[36] = |(datain[167:164] ^ 3);
  assign w954[37] = |(datain[163:160] ^ 12);
  assign w954[38] = |(datain[159:156] ^ 0);
  assign w954[39] = |(datain[155:152] ^ 0);
  assign w954[40] = |(datain[151:148] ^ 7);
  assign w954[41] = |(datain[147:144] ^ 4);
  assign w954[42] = |(datain[143:140] ^ 0);
  assign w954[43] = |(datain[139:136] ^ 5);
  assign w954[44] = |(datain[135:132] ^ 0);
  assign w954[45] = |(datain[131:128] ^ 14);
  assign w954[46] = |(datain[127:124] ^ 1);
  assign w954[47] = |(datain[123:120] ^ 15);
  assign w954[48] = |(datain[119:116] ^ 14);
  assign w954[49] = |(datain[115:112] ^ 8);
  assign w954[50] = |(datain[111:108] ^ 0);
  assign w954[51] = |(datain[107:104] ^ 8);
  assign w954[52] = |(datain[103:100] ^ 0);
  assign w954[53] = |(datain[99:96] ^ 0);
  assign w954[54] = |(datain[95:92] ^ 1);
  assign w954[55] = |(datain[91:88] ^ 15);
  assign w954[56] = |(datain[87:84] ^ 5);
  assign w954[57] = |(datain[83:80] ^ 8);
  assign w954[58] = |(datain[79:76] ^ 9);
  assign w954[59] = |(datain[75:72] ^ 13);
  assign w954[60] = |(datain[71:68] ^ 2);
  assign w954[61] = |(datain[67:64] ^ 14);
  assign w954[62] = |(datain[63:60] ^ 15);
  assign w954[63] = |(datain[59:56] ^ 15);
  assign w954[64] = |(datain[55:52] ^ 2);
  assign w954[65] = |(datain[51:48] ^ 14);
  assign w954[66] = |(datain[47:44] ^ 12);
  assign w954[67] = |(datain[43:40] ^ 5);
  assign w954[68] = |(datain[39:36] ^ 0);
  assign w954[69] = |(datain[35:32] ^ 0);
  assign comp[954] = ~(|w954);
  wire [76-1:0] w955;
  assign w955[0] = |(datain[311:308] ^ 0);
  assign w955[1] = |(datain[307:304] ^ 3);
  assign w955[2] = |(datain[303:300] ^ 11);
  assign w955[3] = |(datain[299:296] ^ 14);
  assign w955[4] = |(datain[295:292] ^ 0);
  assign w955[5] = |(datain[291:288] ^ 0);
  assign w955[6] = |(datain[287:284] ^ 0);
  assign w955[7] = |(datain[283:280] ^ 1);
  assign w955[8] = |(datain[279:276] ^ 11);
  assign w955[9] = |(datain[275:272] ^ 9);
  assign w955[10] = |(datain[271:268] ^ 0);
  assign w955[11] = |(datain[267:264] ^ 6);
  assign w955[12] = |(datain[263:260] ^ 0);
  assign w955[13] = |(datain[259:256] ^ 0);
  assign w955[14] = |(datain[255:252] ^ 15);
  assign w955[15] = |(datain[251:248] ^ 12);
  assign w955[16] = |(datain[247:244] ^ 10);
  assign w955[17] = |(datain[243:240] ^ 6);
  assign w955[18] = |(datain[239:236] ^ 7);
  assign w955[19] = |(datain[235:232] ^ 5);
  assign w955[20] = |(datain[231:228] ^ 0);
  assign w955[21] = |(datain[227:224] ^ 4);
  assign w955[22] = |(datain[223:220] ^ 14);
  assign w955[23] = |(datain[219:216] ^ 2);
  assign w955[24] = |(datain[215:212] ^ 15);
  assign w955[25] = |(datain[211:208] ^ 11);
  assign w955[26] = |(datain[207:204] ^ 14);
  assign w955[27] = |(datain[203:200] ^ 11);
  assign w955[28] = |(datain[199:196] ^ 7);
  assign w955[29] = |(datain[195:192] ^ 0);
  assign w955[30] = |(datain[191:188] ^ 8);
  assign w955[31] = |(datain[187:184] ^ 0);
  assign w955[32] = |(datain[183:180] ^ 15);
  assign w955[33] = |(datain[179:176] ^ 10);
  assign w955[34] = |(datain[175:172] ^ 8);
  assign w955[35] = |(datain[171:168] ^ 0);
  assign w955[36] = |(datain[167:164] ^ 7);
  assign w955[37] = |(datain[163:160] ^ 2);
  assign w955[38] = |(datain[159:156] ^ 1);
  assign w955[39] = |(datain[155:152] ^ 3);
  assign w955[40] = |(datain[151:148] ^ 11);
  assign w955[41] = |(datain[147:144] ^ 6);
  assign w955[42] = |(datain[143:140] ^ 0);
  assign w955[43] = |(datain[139:136] ^ 0);
  assign w955[44] = |(datain[135:132] ^ 11);
  assign w955[45] = |(datain[131:128] ^ 9);
  assign w955[46] = |(datain[127:124] ^ 0);
  assign w955[47] = |(datain[123:120] ^ 6);
  assign w955[48] = |(datain[119:116] ^ 0);
  assign w955[49] = |(datain[115:112] ^ 0);
  assign w955[50] = |(datain[111:108] ^ 11);
  assign w955[51] = |(datain[107:104] ^ 8);
  assign w955[52] = |(datain[103:100] ^ 0);
  assign w955[53] = |(datain[99:96] ^ 1);
  assign w955[54] = |(datain[95:92] ^ 0);
  assign w955[55] = |(datain[91:88] ^ 3);
  assign w955[56] = |(datain[87:84] ^ 5);
  assign w955[57] = |(datain[83:80] ^ 1);
  assign w955[58] = |(datain[79:76] ^ 5);
  assign w955[59] = |(datain[75:72] ^ 2);
  assign w955[60] = |(datain[71:68] ^ 9);
  assign w955[61] = |(datain[67:64] ^ 12);
  assign w955[62] = |(datain[63:60] ^ 15);
  assign w955[63] = |(datain[59:56] ^ 15);
  assign w955[64] = |(datain[55:52] ^ 1);
  assign w955[65] = |(datain[51:48] ^ 14);
  assign w955[66] = |(datain[47:44] ^ 12);
  assign w955[67] = |(datain[43:40] ^ 5);
  assign w955[68] = |(datain[39:36] ^ 0);
  assign w955[69] = |(datain[35:32] ^ 0);
  assign w955[70] = |(datain[31:28] ^ 7);
  assign w955[71] = |(datain[27:24] ^ 3);
  assign w955[72] = |(datain[23:20] ^ 3);
  assign w955[73] = |(datain[19:16] ^ 1);
  assign w955[74] = |(datain[15:12] ^ 14);
  assign w955[75] = |(datain[11:8] ^ 11);
  assign comp[955] = ~(|w955);
  wire [76-1:0] w956;
  assign w956[0] = |(datain[311:308] ^ 11);
  assign w956[1] = |(datain[307:304] ^ 15);
  assign w956[2] = |(datain[303:300] ^ 7);
  assign w956[3] = |(datain[299:296] ^ 12);
  assign w956[4] = |(datain[295:292] ^ 3);
  assign w956[5] = |(datain[291:288] ^ 3);
  assign w956[6] = |(datain[287:284] ^ 12);
  assign w956[7] = |(datain[283:280] ^ 0);
  assign w956[8] = |(datain[279:276] ^ 12);
  assign w956[9] = |(datain[275:272] ^ 13);
  assign w956[10] = |(datain[271:268] ^ 1);
  assign w956[11] = |(datain[267:264] ^ 3);
  assign w956[12] = |(datain[263:260] ^ 8);
  assign w956[13] = |(datain[259:256] ^ 14);
  assign w956[14] = |(datain[255:252] ^ 12);
  assign w956[15] = |(datain[251:248] ^ 0);
  assign w956[16] = |(datain[247:244] ^ 0);
  assign w956[17] = |(datain[243:240] ^ 14);
  assign w956[18] = |(datain[239:236] ^ 1);
  assign w956[19] = |(datain[235:232] ^ 15);
  assign w956[20] = |(datain[231:228] ^ 11);
  assign w956[21] = |(datain[227:224] ^ 11);
  assign w956[22] = |(datain[223:220] ^ 0);
  assign w956[23] = |(datain[219:216] ^ 0);
  assign w956[24] = |(datain[215:212] ^ 7);
  assign w956[25] = |(datain[211:208] ^ 12);
  assign w956[26] = |(datain[207:204] ^ 11);
  assign w956[27] = |(datain[203:200] ^ 8);
  assign w956[28] = |(datain[199:196] ^ 0);
  assign w956[29] = |(datain[195:192] ^ 1);
  assign w956[30] = |(datain[191:188] ^ 0);
  assign w956[31] = |(datain[187:184] ^ 2);
  assign w956[32] = |(datain[183:180] ^ 11);
  assign w956[33] = |(datain[179:176] ^ 5);
  assign w956[34] = |(datain[175:172] ^ 0);
  assign w956[35] = |(datain[171:168] ^ 0);
  assign w956[36] = |(datain[167:164] ^ 8);
  assign w956[37] = |(datain[163:160] ^ 0);
  assign w956[38] = |(datain[159:156] ^ 3);
  assign w956[39] = |(datain[155:152] ^ 14);
  assign w956[40] = |(datain[151:148] ^ 12);
  assign w956[41] = |(datain[147:144] ^ 3);
  assign w956[42] = |(datain[143:140] ^ 0);
  assign w956[43] = |(datain[139:136] ^ 0);
  assign w956[44] = |(datain[135:132] ^ 8);
  assign w956[45] = |(datain[131:128] ^ 0);
  assign w956[46] = |(datain[127:124] ^ 9);
  assign w956[47] = |(datain[123:120] ^ 0);
  assign w956[48] = |(datain[119:116] ^ 7);
  assign w956[49] = |(datain[115:112] ^ 3);
  assign w956[50] = |(datain[111:108] ^ 1);
  assign w956[51] = |(datain[107:104] ^ 7);
  assign w956[52] = |(datain[103:100] ^ 11);
  assign w956[53] = |(datain[99:96] ^ 6);
  assign w956[54] = |(datain[95:92] ^ 0);
  assign w956[55] = |(datain[91:88] ^ 1);
  assign w956[56] = |(datain[87:84] ^ 8);
  assign w956[57] = |(datain[83:80] ^ 10);
  assign w956[58] = |(datain[79:76] ^ 1);
  assign w956[59] = |(datain[75:72] ^ 6);
  assign w956[60] = |(datain[71:68] ^ 12);
  assign w956[61] = |(datain[67:64] ^ 3);
  assign w956[62] = |(datain[63:60] ^ 0);
  assign w956[63] = |(datain[59:56] ^ 0);
  assign w956[64] = |(datain[55:52] ^ 8);
  assign w956[65] = |(datain[51:48] ^ 10);
  assign w956[66] = |(datain[47:44] ^ 0);
  assign w956[67] = |(datain[43:40] ^ 14);
  assign w956[68] = |(datain[39:36] ^ 12);
  assign w956[69] = |(datain[35:32] ^ 4);
  assign w956[70] = |(datain[31:28] ^ 0);
  assign w956[71] = |(datain[27:24] ^ 0);
  assign w956[72] = |(datain[23:20] ^ 12);
  assign w956[73] = |(datain[19:16] ^ 13);
  assign w956[74] = |(datain[15:12] ^ 1);
  assign w956[75] = |(datain[11:8] ^ 3);
  assign comp[956] = ~(|w956);
  wire [32-1:0] w957;
  assign w957[0] = |(datain[311:308] ^ 11);
  assign w957[1] = |(datain[307:304] ^ 11);
  assign w957[2] = |(datain[303:300] ^ 1);
  assign w957[3] = |(datain[299:296] ^ 0);
  assign w957[4] = |(datain[295:292] ^ 0);
  assign w957[5] = |(datain[291:288] ^ 0);
  assign w957[6] = |(datain[287:284] ^ 11);
  assign w957[7] = |(datain[283:280] ^ 9);
  assign w957[8] = |(datain[279:276] ^ 14);
  assign w957[9] = |(datain[275:272] ^ 8);
  assign w957[10] = |(datain[271:268] ^ 0);
  assign w957[11] = |(datain[267:264] ^ 3);
  assign w957[12] = |(datain[263:260] ^ 11);
  assign w957[13] = |(datain[259:256] ^ 0);
  assign w957[14] = |(datain[255:252] ^ 15);
  assign w957[15] = |(datain[251:248] ^ 12);
  assign w957[16] = |(datain[247:244] ^ 2);
  assign w957[17] = |(datain[243:240] ^ 14);
  assign w957[18] = |(datain[239:236] ^ 0);
  assign w957[19] = |(datain[235:232] ^ 0);
  assign w957[20] = |(datain[231:228] ^ 0);
  assign w957[21] = |(datain[227:224] ^ 7);
  assign w957[22] = |(datain[223:220] ^ 2);
  assign w957[23] = |(datain[219:216] ^ 10);
  assign w957[24] = |(datain[215:212] ^ 12);
  assign w957[25] = |(datain[211:208] ^ 1);
  assign w957[26] = |(datain[207:204] ^ 4);
  assign w957[27] = |(datain[203:200] ^ 3);
  assign w957[28] = |(datain[199:196] ^ 14);
  assign w957[29] = |(datain[195:192] ^ 2);
  assign w957[30] = |(datain[191:188] ^ 15);
  assign w957[31] = |(datain[187:184] ^ 8);
  assign comp[957] = ~(|w957);
  wire [74-1:0] w958;
  assign w958[0] = |(datain[311:308] ^ 2);
  assign w958[1] = |(datain[307:304] ^ 13);
  assign w958[2] = |(datain[303:300] ^ 0);
  assign w958[3] = |(datain[299:296] ^ 2);
  assign w958[4] = |(datain[295:292] ^ 0);
  assign w958[5] = |(datain[291:288] ^ 0);
  assign w958[6] = |(datain[287:284] ^ 10);
  assign w958[7] = |(datain[283:280] ^ 3);
  assign w958[8] = |(datain[279:276] ^ 1);
  assign w958[9] = |(datain[275:272] ^ 3);
  assign w958[10] = |(datain[271:268] ^ 0);
  assign w958[11] = |(datain[267:264] ^ 4);
  assign w958[12] = |(datain[263:260] ^ 11);
  assign w958[13] = |(datain[259:256] ^ 1);
  assign w958[14] = |(datain[255:252] ^ 0);
  assign w958[15] = |(datain[251:248] ^ 6);
  assign w958[16] = |(datain[247:244] ^ 13);
  assign w958[17] = |(datain[243:240] ^ 3);
  assign w958[18] = |(datain[239:236] ^ 14);
  assign w958[19] = |(datain[235:232] ^ 0);
  assign w958[20] = |(datain[231:228] ^ 2);
  assign w958[21] = |(datain[227:224] ^ 13);
  assign w958[22] = |(datain[223:220] ^ 6);
  assign w958[23] = |(datain[219:216] ^ 0);
  assign w958[24] = |(datain[215:212] ^ 0);
  assign w958[25] = |(datain[211:208] ^ 0);
  assign w958[26] = |(datain[207:204] ^ 8);
  assign w958[27] = |(datain[203:200] ^ 14);
  assign w958[28] = |(datain[199:196] ^ 12);
  assign w958[29] = |(datain[195:192] ^ 0);
  assign w958[30] = |(datain[191:188] ^ 8);
  assign w958[31] = |(datain[187:184] ^ 11);
  assign w958[32] = |(datain[183:180] ^ 15);
  assign w958[33] = |(datain[179:176] ^ 4);
  assign w958[34] = |(datain[175:172] ^ 11);
  assign w958[35] = |(datain[171:168] ^ 15);
  assign w958[36] = |(datain[167:164] ^ 0);
  assign w958[37] = |(datain[163:160] ^ 4);
  assign w958[38] = |(datain[159:156] ^ 0);
  assign w958[39] = |(datain[155:152] ^ 6);
  assign w958[40] = |(datain[151:148] ^ 11);
  assign w958[41] = |(datain[147:144] ^ 9);
  assign w958[42] = |(datain[143:140] ^ 0);
  assign w958[43] = |(datain[139:136] ^ 0);
  assign w958[44] = |(datain[135:132] ^ 0);
  assign w958[45] = |(datain[131:128] ^ 1);
  assign w958[46] = |(datain[127:124] ^ 15);
  assign w958[47] = |(datain[123:120] ^ 3);
  assign w958[48] = |(datain[119:116] ^ 10);
  assign w958[49] = |(datain[115:112] ^ 5);
  assign w958[50] = |(datain[111:108] ^ 11);
  assign w958[51] = |(datain[107:104] ^ 10);
  assign w958[52] = |(datain[103:100] ^ 7);
  assign w958[53] = |(datain[99:96] ^ 11);
  assign w958[54] = |(datain[95:92] ^ 0);
  assign w958[55] = |(datain[91:88] ^ 6);
  assign w958[56] = |(datain[87:84] ^ 0);
  assign w958[57] = |(datain[83:80] ^ 6);
  assign w958[58] = |(datain[79:76] ^ 5);
  assign w958[59] = |(datain[75:72] ^ 2);
  assign w958[60] = |(datain[71:68] ^ 12);
  assign w958[61] = |(datain[67:64] ^ 11);
  assign w958[62] = |(datain[63:60] ^ 3);
  assign w958[63] = |(datain[59:56] ^ 3);
  assign w958[64] = |(datain[55:52] ^ 12);
  assign w958[65] = |(datain[51:48] ^ 0);
  assign w958[66] = |(datain[47:44] ^ 2);
  assign w958[67] = |(datain[43:40] ^ 2);
  assign w958[68] = |(datain[39:36] ^ 13);
  assign w958[69] = |(datain[35:32] ^ 0);
  assign w958[70] = |(datain[31:28] ^ 12);
  assign w958[71] = |(datain[27:24] ^ 13);
  assign w958[72] = |(datain[23:20] ^ 1);
  assign w958[73] = |(datain[19:16] ^ 3);
  assign comp[958] = ~(|w958);
  wire [76-1:0] w959;
  assign w959[0] = |(datain[311:308] ^ 0);
  assign w959[1] = |(datain[307:304] ^ 4);
  assign w959[2] = |(datain[303:300] ^ 8);
  assign w959[3] = |(datain[299:296] ^ 3);
  assign w959[4] = |(datain[295:292] ^ 4);
  assign w959[5] = |(datain[291:288] ^ 4);
  assign w959[6] = |(datain[287:284] ^ 0);
  assign w959[7] = |(datain[283:280] ^ 1);
  assign w959[8] = |(datain[279:276] ^ 15);
  assign w959[9] = |(datain[275:272] ^ 13);
  assign w959[10] = |(datain[271:268] ^ 10);
  assign w959[11] = |(datain[267:264] ^ 12);
  assign w959[12] = |(datain[263:260] ^ 10);
  assign w959[13] = |(datain[259:256] ^ 13);
  assign w959[14] = |(datain[255:252] ^ 11);
  assign w959[15] = |(datain[251:248] ^ 1);
  assign w959[16] = |(datain[247:244] ^ 0);
  assign w959[17] = |(datain[243:240] ^ 6);
  assign w959[18] = |(datain[239:236] ^ 13);
  assign w959[19] = |(datain[235:232] ^ 3);
  assign w959[20] = |(datain[231:228] ^ 14);
  assign w959[21] = |(datain[227:224] ^ 0);
  assign w959[22] = |(datain[223:220] ^ 8);
  assign w959[23] = |(datain[219:216] ^ 14);
  assign w959[24] = |(datain[215:212] ^ 12);
  assign w959[25] = |(datain[211:208] ^ 0);
  assign w959[26] = |(datain[207:204] ^ 3);
  assign w959[27] = |(datain[203:200] ^ 3);
  assign w959[28] = |(datain[199:196] ^ 13);
  assign w959[29] = |(datain[195:192] ^ 11);
  assign w959[30] = |(datain[191:188] ^ 11);
  assign w959[31] = |(datain[187:184] ^ 8);
  assign w959[32] = |(datain[183:180] ^ 0);
  assign w959[33] = |(datain[179:176] ^ 4);
  assign w959[34] = |(datain[175:172] ^ 0);
  assign w959[35] = |(datain[171:168] ^ 2);
  assign w959[36] = |(datain[167:164] ^ 5);
  assign w959[37] = |(datain[163:160] ^ 9);
  assign w959[38] = |(datain[159:156] ^ 5);
  assign w959[39] = |(datain[155:152] ^ 1);
  assign w959[40] = |(datain[151:148] ^ 4);
  assign w959[41] = |(datain[147:144] ^ 1);
  assign w959[42] = |(datain[143:140] ^ 12);
  assign w959[43] = |(datain[139:136] ^ 13);
  assign w959[44] = |(datain[135:132] ^ 1);
  assign w959[45] = |(datain[131:128] ^ 3);
  assign w959[46] = |(datain[127:124] ^ 0);
  assign w959[47] = |(datain[123:120] ^ 6);
  assign w959[48] = |(datain[119:116] ^ 11);
  assign w959[49] = |(datain[115:112] ^ 8);
  assign w959[50] = |(datain[111:108] ^ 5);
  assign w959[51] = |(datain[107:104] ^ 7);
  assign w959[52] = |(datain[103:100] ^ 0);
  assign w959[53] = |(datain[99:96] ^ 7);
  assign w959[54] = |(datain[95:92] ^ 5);
  assign w959[55] = |(datain[91:88] ^ 0);
  assign w959[56] = |(datain[87:84] ^ 12);
  assign w959[57] = |(datain[83:80] ^ 11);
  assign w959[58] = |(datain[79:76] ^ 11);
  assign w959[59] = |(datain[75:72] ^ 8);
  assign w959[60] = |(datain[71:68] ^ 12);
  assign w959[61] = |(datain[67:64] ^ 14);
  assign w959[62] = |(datain[63:60] ^ 10);
  assign w959[63] = |(datain[59:56] ^ 7);
  assign w959[64] = |(datain[55:52] ^ 12);
  assign w959[65] = |(datain[51:48] ^ 13);
  assign w959[66] = |(datain[47:44] ^ 1);
  assign w959[67] = |(datain[43:40] ^ 3);
  assign w959[68] = |(datain[39:36] ^ 8);
  assign w959[69] = |(datain[35:32] ^ 1);
  assign w959[70] = |(datain[31:28] ^ 15);
  assign w959[71] = |(datain[27:24] ^ 3);
  assign w959[72] = |(datain[23:20] ^ 12);
  assign w959[73] = |(datain[19:16] ^ 14);
  assign w959[74] = |(datain[15:12] ^ 10);
  assign w959[75] = |(datain[11:8] ^ 7);
  assign comp[959] = ~(|w959);
  wire [46-1:0] w960;
  assign w960[0] = |(datain[311:308] ^ 3);
  assign w960[1] = |(datain[307:304] ^ 3);
  assign w960[2] = |(datain[303:300] ^ 12);
  assign w960[3] = |(datain[299:296] ^ 0);
  assign w960[4] = |(datain[295:292] ^ 8);
  assign w960[5] = |(datain[291:288] ^ 14);
  assign w960[6] = |(datain[287:284] ^ 13);
  assign w960[7] = |(datain[283:280] ^ 8);
  assign w960[8] = |(datain[279:276] ^ 11);
  assign w960[9] = |(datain[275:272] ^ 11);
  assign w960[10] = |(datain[271:268] ^ 2);
  assign w960[11] = |(datain[267:264] ^ 10);
  assign w960[12] = |(datain[263:260] ^ 0);
  assign w960[13] = |(datain[259:256] ^ 1);
  assign w960[14] = |(datain[255:252] ^ 11);
  assign w960[15] = |(datain[251:248] ^ 14);
  assign w960[16] = |(datain[247:244] ^ 0);
  assign w960[17] = |(datain[243:240] ^ 0);
  assign w960[18] = |(datain[239:236] ^ 7);
  assign w960[19] = |(datain[235:232] ^ 12);
  assign w960[20] = |(datain[231:228] ^ 5);
  assign w960[21] = |(datain[227:224] ^ 6);
  assign w960[22] = |(datain[223:220] ^ 15);
  assign w960[23] = |(datain[219:216] ^ 15);
  assign w960[24] = |(datain[215:212] ^ 0);
  assign w960[25] = |(datain[211:208] ^ 14);
  assign w960[26] = |(datain[207:204] ^ 1);
  assign w960[27] = |(datain[203:200] ^ 3);
  assign w960[28] = |(datain[199:196] ^ 0);
  assign w960[29] = |(datain[195:192] ^ 4);
  assign w960[30] = |(datain[191:188] ^ 10);
  assign w960[31] = |(datain[187:184] ^ 1);
  assign w960[32] = |(datain[183:180] ^ 1);
  assign w960[33] = |(datain[179:176] ^ 3);
  assign w960[34] = |(datain[175:172] ^ 0);
  assign w960[35] = |(datain[171:168] ^ 4);
  assign w960[36] = |(datain[167:164] ^ 12);
  assign w960[37] = |(datain[163:160] ^ 1);
  assign w960[38] = |(datain[159:156] ^ 14);
  assign w960[39] = |(datain[155:152] ^ 0);
  assign w960[40] = |(datain[151:148] ^ 0);
  assign w960[41] = |(datain[147:144] ^ 6);
  assign w960[42] = |(datain[143:140] ^ 2);
  assign w960[43] = |(datain[139:136] ^ 13);
  assign w960[44] = |(datain[135:132] ^ 1);
  assign w960[45] = |(datain[131:128] ^ 0);
  assign comp[960] = ~(|w960);
  wire [76-1:0] w961;
  assign w961[0] = |(datain[311:308] ^ 0);
  assign w961[1] = |(datain[307:304] ^ 2);
  assign w961[2] = |(datain[303:300] ^ 11);
  assign w961[3] = |(datain[299:296] ^ 9);
  assign w961[4] = |(datain[295:292] ^ 0);
  assign w961[5] = |(datain[291:288] ^ 1);
  assign w961[6] = |(datain[287:284] ^ 0);
  assign w961[7] = |(datain[283:280] ^ 0);
  assign w961[8] = |(datain[279:276] ^ 11);
  assign w961[9] = |(datain[275:272] ^ 10);
  assign w961[10] = |(datain[271:268] ^ 8);
  assign w961[11] = |(datain[267:264] ^ 0);
  assign w961[12] = |(datain[263:260] ^ 0);
  assign w961[13] = |(datain[259:256] ^ 0);
  assign w961[14] = |(datain[255:252] ^ 12);
  assign w961[15] = |(datain[251:248] ^ 13);
  assign w961[16] = |(datain[247:244] ^ 1);
  assign w961[17] = |(datain[243:240] ^ 3);
  assign w961[18] = |(datain[239:236] ^ 7);
  assign w961[19] = |(datain[235:232] ^ 2);
  assign w961[20] = |(datain[231:228] ^ 1);
  assign w961[21] = |(datain[227:224] ^ 10);
  assign w961[22] = |(datain[223:220] ^ 2);
  assign w961[23] = |(datain[219:216] ^ 6);
  assign w961[24] = |(datain[215:212] ^ 8);
  assign w961[25] = |(datain[211:208] ^ 0);
  assign w961[26] = |(datain[207:204] ^ 3);
  assign w961[27] = |(datain[203:200] ^ 15);
  assign w961[28] = |(datain[199:196] ^ 14);
  assign w961[29] = |(datain[195:192] ^ 8);
  assign w961[30] = |(datain[191:188] ^ 7);
  assign w961[31] = |(datain[187:184] ^ 4);
  assign w961[32] = |(datain[183:180] ^ 1);
  assign w961[33] = |(datain[179:176] ^ 4);
  assign w961[34] = |(datain[175:172] ^ 11);
  assign w961[35] = |(datain[171:168] ^ 8);
  assign w961[36] = |(datain[167:164] ^ 0);
  assign w961[37] = |(datain[163:160] ^ 1);
  assign w961[38] = |(datain[159:156] ^ 0);
  assign w961[39] = |(datain[155:152] ^ 3);
  assign w961[40] = |(datain[151:148] ^ 4);
  assign w961[41] = |(datain[147:144] ^ 1);
  assign w961[42] = |(datain[143:140] ^ 12);
  assign w961[43] = |(datain[139:136] ^ 13);
  assign w961[44] = |(datain[135:132] ^ 1);
  assign w961[45] = |(datain[131:128] ^ 3);
  assign w961[46] = |(datain[127:124] ^ 8);
  assign w961[47] = |(datain[123:120] ^ 9);
  assign w961[48] = |(datain[119:116] ^ 13);
  assign w961[49] = |(datain[115:112] ^ 15);
  assign w961[50] = |(datain[111:108] ^ 11);
  assign w961[51] = |(datain[107:104] ^ 9);
  assign w961[52] = |(datain[103:100] ^ 11);
  assign w961[53] = |(datain[99:96] ^ 10);
  assign w961[54] = |(datain[95:92] ^ 0);
  assign w961[55] = |(datain[91:88] ^ 1);
  assign w961[56] = |(datain[87:84] ^ 15);
  assign w961[57] = |(datain[83:80] ^ 12);
  assign w961[58] = |(datain[79:76] ^ 15);
  assign w961[59] = |(datain[75:72] ^ 3);
  assign w961[60] = |(datain[71:68] ^ 10);
  assign w961[61] = |(datain[67:64] ^ 4);
  assign w961[62] = |(datain[63:60] ^ 11);
  assign w961[63] = |(datain[59:56] ^ 8);
  assign w961[64] = |(datain[55:52] ^ 0);
  assign w961[65] = |(datain[51:48] ^ 1);
  assign w961[66] = |(datain[47:44] ^ 0);
  assign w961[67] = |(datain[43:40] ^ 3);
  assign w961[68] = |(datain[39:36] ^ 4);
  assign w961[69] = |(datain[35:32] ^ 1);
  assign w961[70] = |(datain[31:28] ^ 12);
  assign w961[71] = |(datain[27:24] ^ 13);
  assign w961[72] = |(datain[23:20] ^ 1);
  assign w961[73] = |(datain[19:16] ^ 3);
  assign w961[74] = |(datain[15:12] ^ 11);
  assign w961[75] = |(datain[11:8] ^ 8);
  assign comp[961] = ~(|w961);
  wire [54-1:0] w962;
  assign w962[0] = |(datain[311:308] ^ 12);
  assign w962[1] = |(datain[307:304] ^ 0);
  assign w962[2] = |(datain[303:300] ^ 8);
  assign w962[3] = |(datain[299:296] ^ 14);
  assign w962[4] = |(datain[295:292] ^ 13);
  assign w962[5] = |(datain[291:288] ^ 0);
  assign w962[6] = |(datain[287:284] ^ 11);
  assign w962[7] = |(datain[283:280] ^ 12);
  assign w962[8] = |(datain[279:276] ^ 0);
  assign w962[9] = |(datain[275:272] ^ 0);
  assign w962[10] = |(datain[271:268] ^ 7);
  assign w962[11] = |(datain[267:264] ^ 12);
  assign w962[12] = |(datain[263:260] ^ 15);
  assign w962[13] = |(datain[259:256] ^ 11);
  assign w962[14] = |(datain[255:252] ^ 8);
  assign w962[15] = |(datain[251:248] ^ 14);
  assign w962[16] = |(datain[247:244] ^ 12);
  assign w962[17] = |(datain[243:240] ^ 0);
  assign w962[18] = |(datain[239:236] ^ 11);
  assign w962[19] = |(datain[235:232] ^ 8);
  assign w962[20] = |(datain[231:228] ^ 0);
  assign w962[21] = |(datain[227:224] ^ 1);
  assign w962[22] = |(datain[223:220] ^ 0);
  assign w962[23] = |(datain[219:216] ^ 2);
  assign w962[24] = |(datain[215:212] ^ 11);
  assign w962[25] = |(datain[211:208] ^ 11);
  assign w962[26] = |(datain[207:204] ^ 0);
  assign w962[27] = |(datain[203:200] ^ 0);
  assign w962[28] = |(datain[199:196] ^ 7);
  assign w962[29] = |(datain[195:192] ^ 14);
  assign w962[30] = |(datain[191:188] ^ 11);
  assign w962[31] = |(datain[187:184] ^ 9);
  assign w962[32] = |(datain[183:180] ^ 0);
  assign w962[33] = |(datain[179:176] ^ 14);
  assign w962[34] = |(datain[175:172] ^ 0);
  assign w962[35] = |(datain[171:168] ^ 0);
  assign w962[36] = |(datain[167:164] ^ 11);
  assign w962[37] = |(datain[163:160] ^ 6);
  assign w962[38] = |(datain[159:156] ^ 0);
  assign w962[39] = |(datain[155:152] ^ 1);
  assign w962[40] = |(datain[151:148] ^ 11);
  assign w962[41] = |(datain[147:144] ^ 2);
  assign w962[42] = |(datain[143:140] ^ 0);
  assign w962[43] = |(datain[139:136] ^ 0);
  assign w962[44] = |(datain[135:132] ^ 12);
  assign w962[45] = |(datain[131:128] ^ 13);
  assign w962[46] = |(datain[127:124] ^ 1);
  assign w962[47] = |(datain[123:120] ^ 3);
  assign w962[48] = |(datain[119:116] ^ 0);
  assign w962[49] = |(datain[115:112] ^ 6);
  assign w962[50] = |(datain[111:108] ^ 5);
  assign w962[51] = |(datain[107:104] ^ 3);
  assign w962[52] = |(datain[103:100] ^ 12);
  assign w962[53] = |(datain[99:96] ^ 11);
  assign comp[962] = ~(|w962);
  wire [32-1:0] w963;
  assign w963[0] = |(datain[311:308] ^ 10);
  assign w963[1] = |(datain[307:304] ^ 13);
  assign w963[2] = |(datain[303:300] ^ 9);
  assign w963[3] = |(datain[299:296] ^ 2);
  assign w963[4] = |(datain[295:292] ^ 0);
  assign w963[5] = |(datain[291:288] ^ 10);
  assign w963[6] = |(datain[287:284] ^ 1);
  assign w963[7] = |(datain[283:280] ^ 6);
  assign w963[8] = |(datain[279:276] ^ 5);
  assign w963[9] = |(datain[275:272] ^ 12);
  assign w963[10] = |(datain[271:268] ^ 0);
  assign w963[11] = |(datain[267:264] ^ 0);
  assign w963[12] = |(datain[263:260] ^ 8);
  assign w963[13] = |(datain[259:256] ^ 13);
  assign w963[14] = |(datain[255:252] ^ 3);
  assign w963[15] = |(datain[251:248] ^ 2);
  assign w963[16] = |(datain[247:244] ^ 11);
  assign w963[17] = |(datain[243:240] ^ 8);
  assign w963[18] = |(datain[239:236] ^ 0);
  assign w963[19] = |(datain[235:232] ^ 1);
  assign w963[20] = |(datain[231:228] ^ 0);
  assign w963[21] = |(datain[227:224] ^ 3);
  assign w963[22] = |(datain[223:220] ^ 5);
  assign w963[23] = |(datain[219:216] ^ 6);
  assign w963[24] = |(datain[215:212] ^ 5);
  assign w963[25] = |(datain[211:208] ^ 1);
  assign w963[26] = |(datain[207:204] ^ 5);
  assign w963[27] = |(datain[203:200] ^ 2);
  assign w963[28] = |(datain[199:196] ^ 12);
  assign w963[29] = |(datain[195:192] ^ 13);
  assign w963[30] = |(datain[191:188] ^ 1);
  assign w963[31] = |(datain[187:184] ^ 3);
  assign comp[963] = ~(|w963);
  wire [76-1:0] w964;
  assign w964[0] = |(datain[311:308] ^ 15);
  assign w964[1] = |(datain[307:304] ^ 15);
  assign w964[2] = |(datain[303:300] ^ 0);
  assign w964[3] = |(datain[299:296] ^ 14);
  assign w964[4] = |(datain[295:292] ^ 1);
  assign w964[5] = |(datain[291:288] ^ 3);
  assign w964[6] = |(datain[287:284] ^ 0);
  assign w964[7] = |(datain[283:280] ^ 4);
  assign w964[8] = |(datain[279:276] ^ 12);
  assign w964[9] = |(datain[275:272] ^ 13);
  assign w964[10] = |(datain[271:268] ^ 1);
  assign w964[11] = |(datain[267:264] ^ 2);
  assign w964[12] = |(datain[263:260] ^ 11);
  assign w964[13] = |(datain[259:256] ^ 9);
  assign w964[14] = |(datain[255:252] ^ 0);
  assign w964[15] = |(datain[251:248] ^ 10);
  assign w964[16] = |(datain[247:244] ^ 0);
  assign w964[17] = |(datain[243:240] ^ 1);
  assign w964[18] = |(datain[239:236] ^ 13);
  assign w964[19] = |(datain[235:232] ^ 3);
  assign w964[20] = |(datain[231:228] ^ 12);
  assign w964[21] = |(datain[227:224] ^ 8);
  assign w964[22] = |(datain[223:220] ^ 8);
  assign w964[23] = |(datain[219:216] ^ 14);
  assign w964[24] = |(datain[215:212] ^ 12);
  assign w964[25] = |(datain[211:208] ^ 0);
  assign w964[26] = |(datain[207:204] ^ 3);
  assign w964[27] = |(datain[203:200] ^ 3);
  assign w964[28] = |(datain[199:196] ^ 15);
  assign w964[29] = |(datain[195:192] ^ 15);
  assign w964[30] = |(datain[191:188] ^ 11);
  assign w964[31] = |(datain[187:184] ^ 14);
  assign w964[32] = |(datain[183:180] ^ 4);
  assign w964[33] = |(datain[179:176] ^ 1);
  assign w964[34] = |(datain[175:172] ^ 7);
  assign w964[35] = |(datain[171:168] ^ 12);
  assign w964[36] = |(datain[167:164] ^ 15);
  assign w964[37] = |(datain[163:160] ^ 12);
  assign w964[38] = |(datain[159:156] ^ 15);
  assign w964[39] = |(datain[155:152] ^ 3);
  assign w964[40] = |(datain[151:148] ^ 10);
  assign w964[41] = |(datain[147:144] ^ 5);
  assign w964[42] = |(datain[143:140] ^ 14);
  assign w964[43] = |(datain[139:136] ^ 8);
  assign w964[44] = |(datain[135:132] ^ 4);
  assign w964[45] = |(datain[131:128] ^ 5);
  assign w964[46] = |(datain[127:124] ^ 0);
  assign w964[47] = |(datain[123:120] ^ 1);
  assign w964[48] = |(datain[119:116] ^ 12);
  assign w964[49] = |(datain[115:112] ^ 13);
  assign w964[50] = |(datain[111:108] ^ 1);
  assign w964[51] = |(datain[107:104] ^ 9);
  assign w964[52] = |(datain[103:100] ^ 11);
  assign w964[53] = |(datain[99:96] ^ 4);
  assign w964[54] = |(datain[95:92] ^ 4);
  assign w964[55] = |(datain[91:88] ^ 10);
  assign w964[56] = |(datain[87:84] ^ 11);
  assign w964[57] = |(datain[83:80] ^ 11);
  assign w964[58] = |(datain[79:76] ^ 2);
  assign w964[59] = |(datain[75:72] ^ 9);
  assign w964[60] = |(datain[71:68] ^ 0);
  assign w964[61] = |(datain[67:64] ^ 0);
  assign w964[62] = |(datain[63:60] ^ 12);
  assign w964[63] = |(datain[59:56] ^ 13);
  assign w964[64] = |(datain[55:52] ^ 2);
  assign w964[65] = |(datain[51:48] ^ 1);
  assign w964[66] = |(datain[47:44] ^ 3);
  assign w964[67] = |(datain[43:40] ^ 3);
  assign w964[68] = |(datain[39:36] ^ 15);
  assign w964[69] = |(datain[35:32] ^ 6);
  assign w964[70] = |(datain[31:28] ^ 15);
  assign w964[71] = |(datain[27:24] ^ 15);
  assign w964[72] = |(datain[23:20] ^ 7);
  assign w964[73] = |(datain[19:16] ^ 4);
  assign w964[74] = |(datain[15:12] ^ 2);
  assign w964[75] = |(datain[11:8] ^ 12);
  assign comp[964] = ~(|w964);
  wire [76-1:0] w965;
  assign w965[0] = |(datain[311:308] ^ 0);
  assign w965[1] = |(datain[307:304] ^ 1);
  assign w965[2] = |(datain[303:300] ^ 11);
  assign w965[3] = |(datain[299:296] ^ 8);
  assign w965[4] = |(datain[295:292] ^ 0);
  assign w965[5] = |(datain[291:288] ^ 1);
  assign w965[6] = |(datain[287:284] ^ 0);
  assign w965[7] = |(datain[283:280] ^ 2);
  assign w965[8] = |(datain[279:276] ^ 12);
  assign w965[9] = |(datain[275:272] ^ 13);
  assign w965[10] = |(datain[271:268] ^ 1);
  assign w965[11] = |(datain[267:264] ^ 3);
  assign w965[12] = |(datain[263:260] ^ 7);
  assign w965[13] = |(datain[259:256] ^ 2);
  assign w965[14] = |(datain[255:252] ^ 15);
  assign w965[15] = |(datain[251:248] ^ 0);
  assign w965[16] = |(datain[247:244] ^ 14);
  assign w965[17] = |(datain[243:240] ^ 8);
  assign w965[18] = |(datain[239:236] ^ 13);
  assign w965[19] = |(datain[235:232] ^ 14);
  assign w965[20] = |(datain[231:228] ^ 0);
  assign w965[21] = |(datain[227:224] ^ 0);
  assign w965[22] = |(datain[223:220] ^ 5);
  assign w965[23] = |(datain[219:216] ^ 10);
  assign w965[24] = |(datain[215:212] ^ 12);
  assign w965[25] = |(datain[211:208] ^ 11);
  assign w965[26] = |(datain[207:204] ^ 11);
  assign w965[27] = |(datain[203:200] ^ 4);
  assign w965[28] = |(datain[199:196] ^ 15);
  assign w965[29] = |(datain[195:192] ^ 0);
  assign w965[30] = |(datain[191:188] ^ 12);
  assign w965[31] = |(datain[187:184] ^ 13);
  assign w965[32] = |(datain[183:180] ^ 1);
  assign w965[33] = |(datain[179:176] ^ 3);
  assign w965[34] = |(datain[175:172] ^ 8);
  assign w965[35] = |(datain[171:168] ^ 0);
  assign w965[36] = |(datain[167:164] ^ 15);
  assign w965[37] = |(datain[163:160] ^ 12);
  assign w965[38] = |(datain[159:156] ^ 1);
  assign w965[39] = |(datain[155:152] ^ 9);
  assign w965[40] = |(datain[151:148] ^ 7);
  assign w965[41] = |(datain[147:144] ^ 4);
  assign w965[42] = |(datain[143:140] ^ 1);
  assign w965[43] = |(datain[139:136] ^ 0);
  assign w965[44] = |(datain[135:132] ^ 8);
  assign w965[45] = |(datain[131:128] ^ 12);
  assign w965[46] = |(datain[127:124] ^ 13);
  assign w965[47] = |(datain[123:120] ^ 8);
  assign w965[48] = |(datain[119:116] ^ 4);
  assign w965[49] = |(datain[115:112] ^ 8);
  assign w965[50] = |(datain[111:108] ^ 8);
  assign w965[51] = |(datain[107:104] ^ 14);
  assign w965[52] = |(datain[103:100] ^ 13);
  assign w965[53] = |(datain[99:96] ^ 8);
  assign w965[54] = |(datain[95:92] ^ 2);
  assign w965[55] = |(datain[91:88] ^ 9);
  assign w965[56] = |(datain[87:84] ^ 1);
  assign w965[57] = |(datain[83:80] ^ 6);
  assign w965[58] = |(datain[79:76] ^ 0);
  assign w965[59] = |(datain[75:72] ^ 3);
  assign w965[60] = |(datain[71:68] ^ 0);
  assign w965[61] = |(datain[67:64] ^ 0);
  assign w965[62] = |(datain[63:60] ^ 2);
  assign w965[63] = |(datain[59:56] ^ 9);
  assign w965[64] = |(datain[55:52] ^ 1);
  assign w965[65] = |(datain[51:48] ^ 6);
  assign w965[66] = |(datain[47:44] ^ 1);
  assign w965[67] = |(datain[43:40] ^ 2);
  assign w965[68] = |(datain[39:36] ^ 0);
  assign w965[69] = |(datain[35:32] ^ 0);
  assign w965[70] = |(datain[31:28] ^ 14);
  assign w965[71] = |(datain[27:24] ^ 8);
  assign w965[72] = |(datain[23:20] ^ 12);
  assign w965[73] = |(datain[19:16] ^ 3);
  assign w965[74] = |(datain[15:12] ^ 0);
  assign w965[75] = |(datain[11:8] ^ 0);
  assign comp[965] = ~(|w965);
  wire [74-1:0] w966;
  assign w966[0] = |(datain[311:308] ^ 1);
  assign w966[1] = |(datain[307:304] ^ 4);
  assign w966[2] = |(datain[303:300] ^ 8);
  assign w966[3] = |(datain[299:296] ^ 11);
  assign w966[4] = |(datain[295:292] ^ 4);
  assign w966[5] = |(datain[291:288] ^ 12);
  assign w966[6] = |(datain[287:284] ^ 0);
  assign w966[7] = |(datain[283:280] ^ 2);
  assign w966[8] = |(datain[279:276] ^ 11);
  assign w966[9] = |(datain[275:272] ^ 8);
  assign w966[10] = |(datain[271:268] ^ 0);
  assign w966[11] = |(datain[267:264] ^ 1);
  assign w966[12] = |(datain[263:260] ^ 0);
  assign w966[13] = |(datain[259:256] ^ 2);
  assign w966[14] = |(datain[255:252] ^ 14);
  assign w966[15] = |(datain[251:248] ^ 8);
  assign w966[16] = |(datain[247:244] ^ 4);
  assign w966[17] = |(datain[243:240] ^ 10);
  assign w966[18] = |(datain[239:236] ^ 0);
  assign w966[19] = |(datain[235:232] ^ 0);
  assign w966[20] = |(datain[231:228] ^ 7);
  assign w966[21] = |(datain[227:224] ^ 2);
  assign w966[22] = |(datain[223:220] ^ 15);
  assign w966[23] = |(datain[219:216] ^ 3);
  assign w966[24] = |(datain[215:212] ^ 14);
  assign w966[25] = |(datain[211:208] ^ 10);
  assign w966[26] = |(datain[207:204] ^ 0);
  assign w966[27] = |(datain[203:200] ^ 0);
  assign w966[28] = |(datain[199:196] ^ 7);
  assign w966[29] = |(datain[195:192] ^ 12);
  assign w966[30] = |(datain[191:188] ^ 0);
  assign w966[31] = |(datain[187:184] ^ 0);
  assign w966[32] = |(datain[183:180] ^ 0);
  assign w966[33] = |(datain[179:176] ^ 0);
  assign w966[34] = |(datain[175:172] ^ 0);
  assign w966[35] = |(datain[171:168] ^ 14);
  assign w966[36] = |(datain[167:164] ^ 11);
  assign w966[37] = |(datain[163:160] ^ 4);
  assign w966[38] = |(datain[159:156] ^ 1);
  assign w966[39] = |(datain[155:152] ^ 3);
  assign w966[40] = |(datain[151:148] ^ 12);
  assign w966[41] = |(datain[147:144] ^ 13);
  assign w966[42] = |(datain[143:140] ^ 2);
  assign w966[43] = |(datain[139:136] ^ 15);
  assign w966[44] = |(datain[135:132] ^ 1);
  assign w966[45] = |(datain[131:128] ^ 15);
  assign w966[46] = |(datain[127:124] ^ 8);
  assign w966[47] = |(datain[123:120] ^ 12);
  assign w966[48] = |(datain[119:116] ^ 0);
  assign w966[49] = |(datain[115:112] ^ 6);
  assign w966[50] = |(datain[111:108] ^ 3);
  assign w966[51] = |(datain[107:104] ^ 8);
  assign w966[52] = |(datain[103:100] ^ 0);
  assign w966[53] = |(datain[99:96] ^ 1);
  assign w966[54] = |(datain[95:92] ^ 8);
  assign w966[55] = |(datain[91:88] ^ 9);
  assign w966[56] = |(datain[87:84] ^ 1);
  assign w966[57] = |(datain[83:80] ^ 14);
  assign w966[58] = |(datain[79:76] ^ 3);
  assign w966[59] = |(datain[75:72] ^ 6);
  assign w966[60] = |(datain[71:68] ^ 0);
  assign w966[61] = |(datain[67:64] ^ 1);
  assign w966[62] = |(datain[63:60] ^ 0);
  assign w966[63] = |(datain[59:56] ^ 14);
  assign w966[64] = |(datain[55:52] ^ 0);
  assign w966[65] = |(datain[51:48] ^ 7);
  assign w966[66] = |(datain[47:44] ^ 11);
  assign w966[67] = |(datain[43:40] ^ 8);
  assign w966[68] = |(datain[39:36] ^ 0);
  assign w966[69] = |(datain[35:32] ^ 1);
  assign w966[70] = |(datain[31:28] ^ 0);
  assign w966[71] = |(datain[27:24] ^ 2);
  assign w966[72] = |(datain[23:20] ^ 8);
  assign w966[73] = |(datain[19:16] ^ 11);
  assign comp[966] = ~(|w966);
  wire [62-1:0] w967;
  assign w967[0] = |(datain[311:308] ^ 1);
  assign w967[1] = |(datain[307:304] ^ 3);
  assign w967[2] = |(datain[303:300] ^ 12);
  assign w967[3] = |(datain[299:296] ^ 13);
  assign w967[4] = |(datain[295:292] ^ 2);
  assign w967[5] = |(datain[291:288] ^ 15);
  assign w967[6] = |(datain[287:284] ^ 0);
  assign w967[7] = |(datain[283:280] ^ 14);
  assign w967[8] = |(datain[279:276] ^ 1);
  assign w967[9] = |(datain[275:272] ^ 15);
  assign w967[10] = |(datain[271:268] ^ 8);
  assign w967[11] = |(datain[267:264] ^ 9);
  assign w967[12] = |(datain[263:260] ^ 1);
  assign w967[13] = |(datain[259:256] ^ 14);
  assign w967[14] = |(datain[255:252] ^ 4);
  assign w967[15] = |(datain[251:248] ^ 0);
  assign w967[16] = |(datain[247:244] ^ 0);
  assign w967[17] = |(datain[243:240] ^ 1);
  assign w967[18] = |(datain[239:236] ^ 8);
  assign w967[19] = |(datain[235:232] ^ 12);
  assign w967[20] = |(datain[231:228] ^ 0);
  assign w967[21] = |(datain[227:224] ^ 6);
  assign w967[22] = |(datain[223:220] ^ 4);
  assign w967[23] = |(datain[219:216] ^ 2);
  assign w967[24] = |(datain[215:212] ^ 0);
  assign w967[25] = |(datain[211:208] ^ 1);
  assign w967[26] = |(datain[207:204] ^ 0);
  assign w967[27] = |(datain[203:200] ^ 14);
  assign w967[28] = |(datain[199:196] ^ 0);
  assign w967[29] = |(datain[195:192] ^ 7);
  assign w967[30] = |(datain[191:188] ^ 11);
  assign w967[31] = |(datain[187:184] ^ 8);
  assign w967[32] = |(datain[183:180] ^ 0);
  assign w967[33] = |(datain[179:176] ^ 1);
  assign w967[34] = |(datain[175:172] ^ 0);
  assign w967[35] = |(datain[171:168] ^ 2);
  assign w967[36] = |(datain[167:164] ^ 8);
  assign w967[37] = |(datain[163:160] ^ 11);
  assign w967[38] = |(datain[159:156] ^ 13);
  assign w967[39] = |(datain[155:152] ^ 8);
  assign w967[40] = |(datain[151:148] ^ 11);
  assign w967[41] = |(datain[147:144] ^ 9);
  assign w967[42] = |(datain[143:140] ^ 0);
  assign w967[43] = |(datain[139:136] ^ 1);
  assign w967[44] = |(datain[135:132] ^ 0);
  assign w967[45] = |(datain[131:128] ^ 0);
  assign w967[46] = |(datain[127:124] ^ 11);
  assign w967[47] = |(datain[123:120] ^ 10);
  assign w967[48] = |(datain[119:116] ^ 8);
  assign w967[49] = |(datain[115:112] ^ 0);
  assign w967[50] = |(datain[111:108] ^ 0);
  assign w967[51] = |(datain[107:104] ^ 0);
  assign w967[52] = |(datain[103:100] ^ 14);
  assign w967[53] = |(datain[99:96] ^ 8);
  assign w967[54] = |(datain[95:92] ^ 2);
  assign w967[55] = |(datain[91:88] ^ 15);
  assign w967[56] = |(datain[87:84] ^ 0);
  assign w967[57] = |(datain[83:80] ^ 0);
  assign w967[58] = |(datain[79:76] ^ 8);
  assign w967[59] = |(datain[75:72] ^ 11);
  assign w967[60] = |(datain[71:68] ^ 15);
  assign w967[61] = |(datain[67:64] ^ 11);
  assign comp[967] = ~(|w967);
  wire [76-1:0] w968;
  assign w968[0] = |(datain[311:308] ^ 4);
  assign w968[1] = |(datain[307:304] ^ 11);
  assign w968[2] = |(datain[303:300] ^ 7);
  assign w968[3] = |(datain[299:296] ^ 5);
  assign w968[4] = |(datain[295:292] ^ 15);
  assign w968[5] = |(datain[291:288] ^ 1);
  assign w968[6] = |(datain[287:284] ^ 5);
  assign w968[7] = |(datain[283:280] ^ 11);
  assign w968[8] = |(datain[279:276] ^ 5);
  assign w968[9] = |(datain[275:272] ^ 14);
  assign w968[10] = |(datain[271:268] ^ 8);
  assign w968[11] = |(datain[267:264] ^ 11);
  assign w968[12] = |(datain[263:260] ^ 12);
  assign w968[13] = |(datain[259:256] ^ 14);
  assign w968[14] = |(datain[255:252] ^ 8);
  assign w968[15] = |(datain[251:248] ^ 1);
  assign w968[16] = |(datain[247:244] ^ 14);
  assign w968[17] = |(datain[243:240] ^ 9);
  assign w968[18] = |(datain[239:236] ^ 0);
  assign w968[19] = |(datain[235:232] ^ 0);
  assign w968[20] = |(datain[231:228] ^ 0);
  assign w968[21] = |(datain[227:224] ^ 5);
  assign w968[22] = |(datain[223:220] ^ 12);
  assign w968[23] = |(datain[219:216] ^ 1);
  assign w968[24] = |(datain[215:212] ^ 14);
  assign w968[25] = |(datain[211:208] ^ 9);
  assign w968[26] = |(datain[207:204] ^ 0);
  assign w968[27] = |(datain[203:200] ^ 2);
  assign w968[28] = |(datain[199:196] ^ 15);
  assign w968[29] = |(datain[195:192] ^ 13);
  assign w968[30] = |(datain[191:188] ^ 10);
  assign w968[31] = |(datain[187:184] ^ 13);
  assign w968[32] = |(datain[183:180] ^ 5);
  assign w968[33] = |(datain[179:176] ^ 1);
  assign w968[34] = |(datain[175:172] ^ 10);
  assign w968[35] = |(datain[171:168] ^ 13);
  assign w968[36] = |(datain[167:164] ^ 8);
  assign w968[37] = |(datain[163:160] ^ 11);
  assign w968[38] = |(datain[159:156] ^ 12);
  assign w968[39] = |(datain[155:152] ^ 8);
  assign w968[40] = |(datain[151:148] ^ 10);
  assign w968[41] = |(datain[147:144] ^ 13);
  assign w968[42] = |(datain[143:140] ^ 8);
  assign w968[43] = |(datain[139:136] ^ 11);
  assign w968[44] = |(datain[135:132] ^ 13);
  assign w968[45] = |(datain[131:128] ^ 0);
  assign w968[46] = |(datain[127:124] ^ 11);
  assign w968[47] = |(datain[123:120] ^ 2);
  assign w968[48] = |(datain[119:116] ^ 8);
  assign w968[49] = |(datain[115:112] ^ 0);
  assign w968[50] = |(datain[111:108] ^ 11);
  assign w968[51] = |(datain[107:104] ^ 14);
  assign w968[52] = |(datain[103:100] ^ 0);
  assign w968[53] = |(datain[99:96] ^ 4);
  assign w968[54] = |(datain[95:92] ^ 0);
  assign w968[55] = |(datain[91:88] ^ 0);
  assign w968[56] = |(datain[87:84] ^ 11);
  assign w968[57] = |(datain[83:80] ^ 8);
  assign w968[58] = |(datain[79:76] ^ 1);
  assign w968[59] = |(datain[75:72] ^ 0);
  assign w968[60] = |(datain[71:68] ^ 0);
  assign w968[61] = |(datain[67:64] ^ 3);
  assign w968[62] = |(datain[63:60] ^ 12);
  assign w968[63] = |(datain[59:56] ^ 13);
  assign w968[64] = |(datain[55:52] ^ 1);
  assign w968[65] = |(datain[51:48] ^ 3);
  assign w968[66] = |(datain[47:44] ^ 15);
  assign w968[67] = |(datain[43:40] ^ 14);
  assign w968[68] = |(datain[39:36] ^ 12);
  assign w968[69] = |(datain[35:32] ^ 6);
  assign w968[70] = |(datain[31:28] ^ 8);
  assign w968[71] = |(datain[27:24] ^ 0);
  assign w968[72] = |(datain[23:20] ^ 15);
  assign w968[73] = |(datain[19:16] ^ 14);
  assign w968[74] = |(datain[15:12] ^ 1);
  assign w968[75] = |(datain[11:8] ^ 0);
  assign comp[968] = ~(|w968);
  wire [76-1:0] w969;
  assign w969[0] = |(datain[311:308] ^ 14);
  assign w969[1] = |(datain[307:304] ^ 6);
  assign w969[2] = |(datain[303:300] ^ 6);
  assign w969[3] = |(datain[299:296] ^ 1);
  assign w969[4] = |(datain[295:292] ^ 11);
  assign w969[5] = |(datain[291:288] ^ 0);
  assign w969[6] = |(datain[287:284] ^ 0);
  assign w969[7] = |(datain[283:280] ^ 0);
  assign w969[8] = |(datain[279:276] ^ 14);
  assign w969[9] = |(datain[275:272] ^ 6);
  assign w969[10] = |(datain[271:268] ^ 7);
  assign w969[11] = |(datain[267:264] ^ 0);
  assign w969[12] = |(datain[263:260] ^ 5);
  assign w969[13] = |(datain[259:256] ^ 0);
  assign w969[14] = |(datain[255:252] ^ 14);
  assign w969[15] = |(datain[251:248] ^ 4);
  assign w969[16] = |(datain[247:244] ^ 7);
  assign w969[17] = |(datain[243:240] ^ 1);
  assign w969[18] = |(datain[239:236] ^ 8);
  assign w969[19] = |(datain[235:232] ^ 8);
  assign w969[20] = |(datain[231:228] ^ 12);
  assign w969[21] = |(datain[227:224] ^ 4);
  assign w969[22] = |(datain[223:220] ^ 14);
  assign w969[23] = |(datain[219:216] ^ 4);
  assign w969[24] = |(datain[215:212] ^ 7);
  assign w969[25] = |(datain[211:208] ^ 1);
  assign w969[26] = |(datain[207:204] ^ 3);
  assign w969[27] = |(datain[203:200] ^ 8);
  assign w969[28] = |(datain[199:196] ^ 14);
  assign w969[29] = |(datain[195:192] ^ 0);
  assign w969[30] = |(datain[191:188] ^ 7);
  assign w969[31] = |(datain[187:184] ^ 4);
  assign w969[32] = |(datain[183:180] ^ 15);
  assign w969[33] = |(datain[179:176] ^ 10);
  assign w969[34] = |(datain[175:172] ^ 5);
  assign w969[35] = |(datain[171:168] ^ 8);
  assign w969[36] = |(datain[167:164] ^ 14);
  assign w969[37] = |(datain[163:160] ^ 6);
  assign w969[38] = |(datain[159:156] ^ 6);
  assign w969[39] = |(datain[155:152] ^ 1);
  assign w969[40] = |(datain[151:148] ^ 12);
  assign w969[41] = |(datain[147:144] ^ 7);
  assign w969[42] = |(datain[143:140] ^ 0);
  assign w969[43] = |(datain[139:136] ^ 7);
  assign w969[44] = |(datain[135:132] ^ 0);
  assign w969[45] = |(datain[131:128] ^ 0);
  assign w969[46] = |(datain[127:124] ^ 1);
  assign w969[47] = |(datain[123:120] ^ 0);
  assign w969[48] = |(datain[119:116] ^ 15);
  assign w969[49] = |(datain[115:112] ^ 14);
  assign w969[50] = |(datain[111:108] ^ 4);
  assign w969[51] = |(datain[107:104] ^ 15);
  assign w969[52] = |(datain[103:100] ^ 0);
  assign w969[53] = |(datain[99:96] ^ 2);
  assign w969[54] = |(datain[95:92] ^ 7);
  assign w969[55] = |(datain[91:88] ^ 5);
  assign w969[56] = |(datain[87:84] ^ 0);
  assign w969[57] = |(datain[83:80] ^ 13);
  assign w969[58] = |(datain[79:76] ^ 5);
  assign w969[59] = |(datain[75:72] ^ 2);
  assign w969[60] = |(datain[71:68] ^ 11);
  assign w969[61] = |(datain[67:64] ^ 8);
  assign w969[62] = |(datain[63:60] ^ 0);
  assign w969[63] = |(datain[59:56] ^ 4);
  assign w969[64] = |(datain[55:52] ^ 0);
  assign w969[65] = |(datain[51:48] ^ 4);
  assign w969[66] = |(datain[47:44] ^ 11);
  assign w969[67] = |(datain[43:40] ^ 10);
  assign w969[68] = |(datain[39:36] ^ 12);
  assign w969[69] = |(datain[35:32] ^ 4);
  assign w969[70] = |(datain[31:28] ^ 0);
  assign w969[71] = |(datain[27:24] ^ 3);
  assign w969[72] = |(datain[23:20] ^ 14);
  assign w969[73] = |(datain[19:16] ^ 15);
  assign w969[74] = |(datain[15:12] ^ 5);
  assign w969[75] = |(datain[11:8] ^ 10);
  assign comp[969] = ~(|w969);
  wire [74-1:0] w970;
  assign w970[0] = |(datain[311:308] ^ 11);
  assign w970[1] = |(datain[307:304] ^ 14);
  assign w970[2] = |(datain[303:300] ^ 0);
  assign w970[3] = |(datain[299:296] ^ 3);
  assign w970[4] = |(datain[295:292] ^ 0);
  assign w970[5] = |(datain[291:288] ^ 0);
  assign w970[6] = |(datain[287:284] ^ 11);
  assign w970[7] = |(datain[283:280] ^ 8);
  assign w970[8] = |(datain[279:276] ^ 0);
  assign w970[9] = |(datain[275:272] ^ 12);
  assign w970[10] = |(datain[271:268] ^ 0);
  assign w970[11] = |(datain[267:264] ^ 2);
  assign w970[12] = |(datain[263:260] ^ 11);
  assign w970[13] = |(datain[259:256] ^ 1);
  assign w970[14] = |(datain[255:252] ^ 0);
  assign w970[15] = |(datain[251:248] ^ 1);
  assign w970[16] = |(datain[247:244] ^ 12);
  assign w970[17] = |(datain[243:240] ^ 13);
  assign w970[18] = |(datain[239:236] ^ 1);
  assign w970[19] = |(datain[235:232] ^ 3);
  assign w970[20] = |(datain[231:228] ^ 4);
  assign w970[21] = |(datain[227:224] ^ 14);
  assign w970[22] = |(datain[223:220] ^ 7);
  assign w970[23] = |(datain[219:216] ^ 4);
  assign w970[24] = |(datain[215:212] ^ 0);
  assign w970[25] = |(datain[211:208] ^ 14);
  assign w970[26] = |(datain[207:204] ^ 7);
  assign w970[27] = |(datain[203:200] ^ 2);
  assign w970[28] = |(datain[199:196] ^ 15);
  assign w970[29] = |(datain[195:192] ^ 4);
  assign w970[30] = |(datain[191:188] ^ 8);
  assign w970[31] = |(datain[187:184] ^ 11);
  assign w970[32] = |(datain[183:180] ^ 14);
  assign w970[33] = |(datain[179:176] ^ 11);
  assign w970[34] = |(datain[175:172] ^ 8);
  assign w970[35] = |(datain[171:168] ^ 1);
  assign w970[36] = |(datain[167:164] ^ 12);
  assign w970[37] = |(datain[163:160] ^ 3);
  assign w970[38] = |(datain[159:156] ^ 3);
  assign w970[39] = |(datain[155:152] ^ 1);
  assign w970[40] = |(datain[151:148] ^ 1);
  assign w970[41] = |(datain[147:144] ^ 2);
  assign w970[42] = |(datain[143:140] ^ 5);
  assign w970[43] = |(datain[139:136] ^ 2);
  assign w970[44] = |(datain[135:132] ^ 5);
  assign w970[45] = |(datain[131:128] ^ 1);
  assign w970[46] = |(datain[127:124] ^ 15);
  assign w970[47] = |(datain[123:120] ^ 15);
  assign w970[48] = |(datain[119:116] ^ 13);
  assign w970[49] = |(datain[115:112] ^ 3);
  assign w970[50] = |(datain[111:108] ^ 5);
  assign w970[51] = |(datain[107:104] ^ 9);
  assign w970[52] = |(datain[103:100] ^ 5);
  assign w970[53] = |(datain[99:96] ^ 10);
  assign w970[54] = |(datain[95:92] ^ 1);
  assign w970[55] = |(datain[91:88] ^ 6);
  assign w970[56] = |(datain[87:84] ^ 0);
  assign w970[57] = |(datain[83:80] ^ 7);
  assign w970[58] = |(datain[79:76] ^ 11);
  assign w970[59] = |(datain[75:72] ^ 8);
  assign w970[60] = |(datain[71:68] ^ 0);
  assign w970[61] = |(datain[67:64] ^ 1);
  assign w970[62] = |(datain[63:60] ^ 0);
  assign w970[63] = |(datain[59:56] ^ 2);
  assign w970[64] = |(datain[55:52] ^ 11);
  assign w970[65] = |(datain[51:48] ^ 11);
  assign w970[66] = |(datain[47:44] ^ 0);
  assign w970[67] = |(datain[43:40] ^ 0);
  assign w970[68] = |(datain[39:36] ^ 7);
  assign w970[69] = |(datain[35:32] ^ 12);
  assign w970[70] = |(datain[31:28] ^ 11);
  assign w970[71] = |(datain[27:24] ^ 1);
  assign w970[72] = |(datain[23:20] ^ 0);
  assign w970[73] = |(datain[19:16] ^ 13);
  assign comp[970] = ~(|w970);
  wire [72-1:0] w971;
  assign w971[0] = |(datain[311:308] ^ 15);
  assign w971[1] = |(datain[307:304] ^ 11);
  assign w971[2] = |(datain[303:300] ^ 8);
  assign w971[3] = |(datain[299:296] ^ 14);
  assign w971[4] = |(datain[295:292] ^ 13);
  assign w971[5] = |(datain[291:288] ^ 8);
  assign w971[6] = |(datain[287:284] ^ 8);
  assign w971[7] = |(datain[283:280] ^ 3);
  assign w971[8] = |(datain[279:276] ^ 2);
  assign w971[9] = |(datain[275:272] ^ 14);
  assign w971[10] = |(datain[271:268] ^ 1);
  assign w971[11] = |(datain[267:264] ^ 3);
  assign w971[12] = |(datain[263:260] ^ 0);
  assign w971[13] = |(datain[259:256] ^ 4);
  assign w971[14] = |(datain[255:252] ^ 0);
  assign w971[15] = |(datain[251:248] ^ 3);
  assign w971[16] = |(datain[247:244] ^ 12);
  assign w971[17] = |(datain[243:240] ^ 13);
  assign w971[18] = |(datain[239:236] ^ 1);
  assign w971[19] = |(datain[235:232] ^ 2);
  assign w971[20] = |(datain[231:228] ^ 11);
  assign w971[21] = |(datain[227:224] ^ 1);
  assign w971[22] = |(datain[223:220] ^ 0);
  assign w971[23] = |(datain[219:216] ^ 6);
  assign w971[24] = |(datain[215:212] ^ 13);
  assign w971[25] = |(datain[211:208] ^ 3);
  assign w971[26] = |(datain[207:204] ^ 14);
  assign w971[27] = |(datain[203:200] ^ 0);
  assign w971[28] = |(datain[199:196] ^ 2);
  assign w971[29] = |(datain[195:192] ^ 13);
  assign w971[30] = |(datain[191:188] ^ 1);
  assign w971[31] = |(datain[187:184] ^ 0);
  assign w971[32] = |(datain[183:180] ^ 0);
  assign w971[33] = |(datain[179:176] ^ 0);
  assign w971[34] = |(datain[175:172] ^ 8);
  assign w971[35] = |(datain[171:168] ^ 14);
  assign w971[36] = |(datain[167:164] ^ 12);
  assign w971[37] = |(datain[163:160] ^ 0);
  assign w971[38] = |(datain[159:156] ^ 11);
  assign w971[39] = |(datain[155:152] ^ 11);
  assign w971[40] = |(datain[151:148] ^ 0);
  assign w971[41] = |(datain[147:144] ^ 0);
  assign w971[42] = |(datain[143:140] ^ 0);
  assign w971[43] = |(datain[139:136] ^ 1);
  assign w971[44] = |(datain[135:132] ^ 11);
  assign w971[45] = |(datain[131:128] ^ 8);
  assign w971[46] = |(datain[127:124] ^ 0);
  assign w971[47] = |(datain[123:120] ^ 3);
  assign w971[48] = |(datain[119:116] ^ 0);
  assign w971[49] = |(datain[115:112] ^ 2);
  assign w971[50] = |(datain[111:108] ^ 11);
  assign w971[51] = |(datain[107:104] ^ 9);
  assign w971[52] = |(datain[103:100] ^ 0);
  assign w971[53] = |(datain[99:96] ^ 3);
  assign w971[54] = |(datain[95:92] ^ 0);
  assign w971[55] = |(datain[91:88] ^ 0);
  assign w971[56] = |(datain[87:84] ^ 11);
  assign w971[57] = |(datain[83:80] ^ 6);
  assign w971[58] = |(datain[79:76] ^ 0);
  assign w971[59] = |(datain[75:72] ^ 0);
  assign w971[60] = |(datain[71:68] ^ 8);
  assign w971[61] = |(datain[67:64] ^ 0);
  assign w971[62] = |(datain[63:60] ^ 15);
  assign w971[63] = |(datain[59:56] ^ 10);
  assign w971[64] = |(datain[55:52] ^ 8);
  assign w971[65] = |(datain[51:48] ^ 0);
  assign w971[66] = |(datain[47:44] ^ 7);
  assign w971[67] = |(datain[43:40] ^ 4);
  assign w971[68] = |(datain[39:36] ^ 0);
  assign w971[69] = |(datain[35:32] ^ 5);
  assign w971[70] = |(datain[31:28] ^ 11);
  assign w971[71] = |(datain[27:24] ^ 9);
  assign comp[971] = ~(|w971);
  wire [76-1:0] w972;
  assign w972[0] = |(datain[311:308] ^ 5);
  assign w972[1] = |(datain[307:304] ^ 3);
  assign w972[2] = |(datain[303:300] ^ 5);
  assign w972[3] = |(datain[299:296] ^ 1);
  assign w972[4] = |(datain[295:292] ^ 1);
  assign w972[5] = |(datain[291:288] ^ 14);
  assign w972[6] = |(datain[287:284] ^ 5);
  assign w972[7] = |(datain[283:280] ^ 6);
  assign w972[8] = |(datain[279:276] ^ 0);
  assign w972[9] = |(datain[275:272] ^ 14);
  assign w972[10] = |(datain[271:268] ^ 1);
  assign w972[11] = |(datain[267:264] ^ 15);
  assign w972[12] = |(datain[263:260] ^ 11);
  assign w972[13] = |(datain[259:256] ^ 4);
  assign w972[14] = |(datain[255:252] ^ 5);
  assign w972[15] = |(datain[251:248] ^ 5);
  assign w972[16] = |(datain[247:244] ^ 11);
  assign w972[17] = |(datain[243:240] ^ 14);
  assign w972[18] = |(datain[239:236] ^ 0);
  assign w972[19] = |(datain[235:232] ^ 0);
  assign w972[20] = |(datain[231:228] ^ 0);
  assign w972[21] = |(datain[227:224] ^ 0);
  assign w972[22] = |(datain[223:220] ^ 11);
  assign w972[23] = |(datain[219:216] ^ 9);
  assign w972[24] = |(datain[215:212] ^ 0);
  assign w972[25] = |(datain[211:208] ^ 0);
  assign w972[26] = |(datain[207:204] ^ 0);
  assign w972[27] = |(datain[203:200] ^ 2);
  assign w972[28] = |(datain[199:196] ^ 8);
  assign w972[29] = |(datain[195:192] ^ 1);
  assign w972[30] = |(datain[191:188] ^ 15);
  assign w972[31] = |(datain[187:184] ^ 14);
  assign w972[32] = |(datain[183:180] ^ 11);
  assign w972[33] = |(datain[179:176] ^ 1);
  assign w972[34] = |(datain[175:172] ^ 0);
  assign w972[35] = |(datain[171:168] ^ 1);
  assign w972[36] = |(datain[167:164] ^ 7);
  assign w972[37] = |(datain[163:160] ^ 2);
  assign w972[38] = |(datain[159:156] ^ 0);
  assign w972[39] = |(datain[155:152] ^ 3);
  assign w972[40] = |(datain[151:148] ^ 11);
  assign w972[41] = |(datain[147:144] ^ 14);
  assign w972[42] = |(datain[143:140] ^ 0);
  assign w972[43] = |(datain[139:136] ^ 0);
  assign w972[44] = |(datain[135:132] ^ 0);
  assign w972[45] = |(datain[131:128] ^ 0);
  assign w972[46] = |(datain[127:124] ^ 3);
  assign w972[47] = |(datain[123:120] ^ 2);
  assign w972[48] = |(datain[119:116] ^ 2);
  assign w972[49] = |(datain[115:112] ^ 4);
  assign w972[50] = |(datain[111:108] ^ 2);
  assign w972[51] = |(datain[107:104] ^ 6);
  assign w972[52] = |(datain[103:100] ^ 3);
  assign w972[53] = |(datain[99:96] ^ 0);
  assign w972[54] = |(datain[95:92] ^ 2);
  assign w972[55] = |(datain[91:88] ^ 7);
  assign w972[56] = |(datain[87:84] ^ 4);
  assign w972[57] = |(datain[83:80] ^ 6);
  assign w972[58] = |(datain[79:76] ^ 4);
  assign w972[59] = |(datain[75:72] ^ 3);
  assign w972[60] = |(datain[71:68] ^ 14);
  assign w972[61] = |(datain[67:64] ^ 2);
  assign w972[62] = |(datain[63:60] ^ 14);
  assign w972[63] = |(datain[59:56] ^ 14);
  assign w972[64] = |(datain[55:52] ^ 15);
  assign w972[65] = |(datain[51:48] ^ 14);
  assign w972[66] = |(datain[47:44] ^ 12);
  assign w972[67] = |(datain[43:40] ^ 8);
  assign w972[68] = |(datain[39:36] ^ 7);
  assign w972[69] = |(datain[35:32] ^ 5);
  assign w972[70] = |(datain[31:28] ^ 14);
  assign w972[71] = |(datain[27:24] ^ 2);
  assign w972[72] = |(datain[23:20] ^ 5);
  assign w972[73] = |(datain[19:16] ^ 14);
  assign w972[74] = |(datain[15:12] ^ 1);
  assign w972[75] = |(datain[11:8] ^ 15);
  assign comp[972] = ~(|w972);
  wire [74-1:0] w973;
  assign w973[0] = |(datain[311:308] ^ 4);
  assign w973[1] = |(datain[307:304] ^ 1);
  assign w973[2] = |(datain[303:300] ^ 14);
  assign w973[3] = |(datain[299:296] ^ 8);
  assign w973[4] = |(datain[295:292] ^ 1);
  assign w973[5] = |(datain[291:288] ^ 5);
  assign w973[6] = |(datain[287:284] ^ 0);
  assign w973[7] = |(datain[283:280] ^ 0);
  assign w973[8] = |(datain[279:276] ^ 5);
  assign w973[9] = |(datain[275:272] ^ 0);
  assign w973[10] = |(datain[271:268] ^ 5);
  assign w973[11] = |(datain[267:264] ^ 0);
  assign w973[12] = |(datain[263:260] ^ 8);
  assign w973[13] = |(datain[259:256] ^ 13);
  assign w973[14] = |(datain[255:252] ^ 11);
  assign w973[15] = |(datain[251:248] ^ 4);
  assign w973[16] = |(datain[247:244] ^ 10);
  assign w973[17] = |(datain[243:240] ^ 15);
  assign w973[18] = |(datain[239:236] ^ 0);
  assign w973[19] = |(datain[235:232] ^ 2);
  assign w973[20] = |(datain[231:228] ^ 11);
  assign w973[21] = |(datain[227:224] ^ 15);
  assign w973[22] = |(datain[223:220] ^ 0);
  assign w973[23] = |(datain[219:216] ^ 0);
  assign w973[24] = |(datain[215:212] ^ 0);
  assign w973[25] = |(datain[211:208] ^ 1);
  assign w973[26] = |(datain[207:204] ^ 5);
  assign w973[27] = |(datain[203:200] ^ 7);
  assign w973[28] = |(datain[199:196] ^ 6);
  assign w973[29] = |(datain[195:192] ^ 6);
  assign w973[30] = |(datain[191:188] ^ 10);
  assign w973[31] = |(datain[187:184] ^ 5);
  assign w973[32] = |(datain[183:180] ^ 3);
  assign w973[33] = |(datain[179:176] ^ 3);
  assign w973[34] = |(datain[175:172] ^ 12);
  assign w973[35] = |(datain[171:168] ^ 0);
  assign w973[36] = |(datain[167:164] ^ 12);
  assign w973[37] = |(datain[163:160] ^ 3);
  assign w973[38] = |(datain[159:156] ^ 11);
  assign w973[39] = |(datain[155:152] ^ 8);
  assign w973[40] = |(datain[151:148] ^ 0);
  assign w973[41] = |(datain[147:144] ^ 1);
  assign w973[42] = |(datain[143:140] ^ 0);
  assign w973[43] = |(datain[139:136] ^ 2);
  assign w973[44] = |(datain[135:132] ^ 11);
  assign w973[45] = |(datain[131:128] ^ 9);
  assign w973[46] = |(datain[127:124] ^ 0);
  assign w973[47] = |(datain[123:120] ^ 1);
  assign w973[48] = |(datain[119:116] ^ 0);
  assign w973[49] = |(datain[115:112] ^ 0);
  assign w973[50] = |(datain[111:108] ^ 11);
  assign w973[51] = |(datain[107:104] ^ 10);
  assign w973[52] = |(datain[103:100] ^ 8);
  assign w973[53] = |(datain[99:96] ^ 0);
  assign w973[54] = |(datain[95:92] ^ 0);
  assign w973[55] = |(datain[91:88] ^ 0);
  assign w973[56] = |(datain[87:84] ^ 12);
  assign w973[57] = |(datain[83:80] ^ 13);
  assign w973[58] = |(datain[79:76] ^ 1);
  assign w973[59] = |(datain[75:72] ^ 3);
  assign w973[60] = |(datain[71:68] ^ 12);
  assign w973[61] = |(datain[67:64] ^ 3);
  assign w973[62] = |(datain[63:60] ^ 8);
  assign w973[63] = |(datain[59:56] ^ 3);
  assign w973[64] = |(datain[55:52] ^ 14);
  assign w973[65] = |(datain[51:48] ^ 10);
  assign w973[66] = |(datain[47:44] ^ 2);
  assign w973[67] = |(datain[43:40] ^ 1);
  assign w973[68] = |(datain[39:36] ^ 12);
  assign w973[69] = |(datain[35:32] ^ 15);
  assign w973[70] = |(datain[31:28] ^ 14);
  assign w973[71] = |(datain[27:24] ^ 11);
  assign w973[72] = |(datain[23:20] ^ 15);
  assign w973[73] = |(datain[19:16] ^ 10);
  assign comp[973] = ~(|w973);
  wire [76-1:0] w974;
  assign w974[0] = |(datain[311:308] ^ 7);
  assign w974[1] = |(datain[307:304] ^ 12);
  assign w974[2] = |(datain[303:300] ^ 3);
  assign w974[3] = |(datain[299:296] ^ 3);
  assign w974[4] = |(datain[295:292] ^ 15);
  assign w974[5] = |(datain[291:288] ^ 15);
  assign w974[6] = |(datain[287:284] ^ 15);
  assign w974[7] = |(datain[283:280] ^ 10);
  assign w974[8] = |(datain[279:276] ^ 8);
  assign w974[9] = |(datain[275:272] ^ 14);
  assign w974[10] = |(datain[271:268] ^ 13);
  assign w974[11] = |(datain[267:264] ^ 7);
  assign w974[12] = |(datain[263:260] ^ 8);
  assign w974[13] = |(datain[259:256] ^ 11);
  assign w974[14] = |(datain[255:252] ^ 14);
  assign w974[15] = |(datain[251:248] ^ 6);
  assign w974[16] = |(datain[247:244] ^ 15);
  assign w974[17] = |(datain[243:240] ^ 11);
  assign w974[18] = |(datain[239:236] ^ 8);
  assign w974[19] = |(datain[235:232] ^ 14);
  assign w974[20] = |(datain[231:228] ^ 13);
  assign w974[21] = |(datain[227:224] ^ 15);
  assign w974[22] = |(datain[223:220] ^ 12);
  assign w974[23] = |(datain[219:216] ^ 6);
  assign w974[24] = |(datain[215:212] ^ 0);
  assign w974[25] = |(datain[211:208] ^ 6);
  assign w974[26] = |(datain[207:204] ^ 1);
  assign w974[27] = |(datain[203:200] ^ 11);
  assign w974[28] = |(datain[199:196] ^ 7);
  assign w974[29] = |(datain[195:192] ^ 12);
  assign w974[30] = |(datain[191:188] ^ 0);
  assign w974[31] = |(datain[187:184] ^ 2);
  assign w974[32] = |(datain[183:180] ^ 12);
  assign w974[33] = |(datain[179:176] ^ 13);
  assign w974[34] = |(datain[175:172] ^ 1);
  assign w974[35] = |(datain[171:168] ^ 2);
  assign w974[36] = |(datain[167:164] ^ 8);
  assign w974[37] = |(datain[163:160] ^ 11);
  assign w974[38] = |(datain[159:156] ^ 14);
  assign w974[39] = |(datain[155:152] ^ 8);
  assign w974[40] = |(datain[151:148] ^ 2);
  assign w974[41] = |(datain[147:144] ^ 13);
  assign w974[42] = |(datain[143:140] ^ 1);
  assign w974[43] = |(datain[139:136] ^ 4);
  assign w974[44] = |(datain[135:132] ^ 0);
  assign w974[45] = |(datain[131:128] ^ 0);
  assign w974[46] = |(datain[127:124] ^ 10);
  assign w974[47] = |(datain[123:120] ^ 3);
  assign w974[48] = |(datain[119:116] ^ 1);
  assign w974[49] = |(datain[115:112] ^ 3);
  assign w974[50] = |(datain[111:108] ^ 0);
  assign w974[51] = |(datain[107:104] ^ 4);
  assign w974[52] = |(datain[103:100] ^ 11);
  assign w974[53] = |(datain[99:96] ^ 1);
  assign w974[54] = |(datain[95:92] ^ 0);
  assign w974[55] = |(datain[91:88] ^ 6);
  assign w974[56] = |(datain[87:84] ^ 13);
  assign w974[57] = |(datain[83:80] ^ 3);
  assign w974[58] = |(datain[79:76] ^ 14);
  assign w974[59] = |(datain[75:72] ^ 0);
  assign w974[60] = |(datain[71:68] ^ 8);
  assign w974[61] = |(datain[67:64] ^ 14);
  assign w974[62] = |(datain[63:60] ^ 12);
  assign w974[63] = |(datain[59:56] ^ 0);
  assign w974[64] = |(datain[55:52] ^ 11);
  assign w974[65] = |(datain[51:48] ^ 9);
  assign w974[66] = |(datain[47:44] ^ 0);
  assign w974[67] = |(datain[43:40] ^ 0);
  assign w974[68] = |(datain[39:36] ^ 0);
  assign w974[69] = |(datain[35:32] ^ 2);
  assign w974[70] = |(datain[31:28] ^ 5);
  assign w974[71] = |(datain[27:24] ^ 1);
  assign w974[72] = |(datain[23:20] ^ 15);
  assign w974[73] = |(datain[19:16] ^ 12);
  assign w974[74] = |(datain[15:12] ^ 15);
  assign w974[75] = |(datain[11:8] ^ 3);
  assign comp[974] = ~(|w974);
  wire [70-1:0] w975;
  assign w975[0] = |(datain[311:308] ^ 15);
  assign w975[1] = |(datain[307:304] ^ 15);
  assign w975[2] = |(datain[303:300] ^ 15);
  assign w975[3] = |(datain[299:296] ^ 10);
  assign w975[4] = |(datain[295:292] ^ 8);
  assign w975[5] = |(datain[291:288] ^ 14);
  assign w975[6] = |(datain[287:284] ^ 13);
  assign w975[7] = |(datain[283:280] ^ 7);
  assign w975[8] = |(datain[279:276] ^ 11);
  assign w975[9] = |(datain[275:272] ^ 12);
  assign w975[10] = |(datain[271:268] ^ 0);
  assign w975[11] = |(datain[267:264] ^ 0);
  assign w975[12] = |(datain[263:260] ^ 7);
  assign w975[13] = |(datain[259:256] ^ 12);
  assign w975[14] = |(datain[255:252] ^ 15);
  assign w975[15] = |(datain[251:248] ^ 11);
  assign w975[16] = |(datain[247:244] ^ 8);
  assign w975[17] = |(datain[243:240] ^ 11);
  assign w975[18] = |(datain[239:236] ^ 15);
  assign w975[19] = |(datain[235:232] ^ 4);
  assign w975[20] = |(datain[231:228] ^ 5);
  assign w975[21] = |(datain[227:224] ^ 7);
  assign w975[22] = |(datain[223:220] ^ 1);
  assign w975[23] = |(datain[219:216] ^ 15);
  assign w975[24] = |(datain[215:212] ^ 15);
  assign w975[25] = |(datain[211:208] ^ 15);
  assign w975[26] = |(datain[207:204] ^ 0);
  assign w975[27] = |(datain[203:200] ^ 14);
  assign w975[28] = |(datain[199:196] ^ 1);
  assign w975[29] = |(datain[195:192] ^ 3);
  assign w975[30] = |(datain[191:188] ^ 0);
  assign w975[31] = |(datain[187:184] ^ 4);
  assign w975[32] = |(datain[183:180] ^ 12);
  assign w975[33] = |(datain[179:176] ^ 13);
  assign w975[34] = |(datain[175:172] ^ 1);
  assign w975[35] = |(datain[171:168] ^ 2);
  assign w975[36] = |(datain[167:164] ^ 12);
  assign w975[37] = |(datain[163:160] ^ 1);
  assign w975[38] = |(datain[159:156] ^ 14);
  assign w975[39] = |(datain[155:152] ^ 0);
  assign w975[40] = |(datain[151:148] ^ 0);
  assign w975[41] = |(datain[147:144] ^ 6);
  assign w975[42] = |(datain[143:140] ^ 5);
  assign w975[43] = |(datain[139:136] ^ 0);
  assign w975[44] = |(datain[135:132] ^ 0);
  assign w975[45] = |(datain[131:128] ^ 7);
  assign w975[46] = |(datain[127:124] ^ 11);
  assign w975[47] = |(datain[123:120] ^ 9);
  assign w975[48] = |(datain[119:116] ^ 0);
  assign w975[49] = |(datain[115:112] ^ 0);
  assign w975[50] = |(datain[111:108] ^ 0);
  assign w975[51] = |(datain[107:104] ^ 2);
  assign w975[52] = |(datain[103:100] ^ 15);
  assign w975[53] = |(datain[99:96] ^ 12);
  assign w975[54] = |(datain[95:92] ^ 15);
  assign w975[55] = |(datain[91:88] ^ 3);
  assign w975[56] = |(datain[87:84] ^ 10);
  assign w975[57] = |(datain[83:80] ^ 5);
  assign w975[58] = |(datain[79:76] ^ 0);
  assign w975[59] = |(datain[75:72] ^ 6);
  assign w975[60] = |(datain[71:68] ^ 11);
  assign w975[61] = |(datain[67:64] ^ 8);
  assign w975[62] = |(datain[63:60] ^ 6);
  assign w975[63] = |(datain[59:56] ^ 2);
  assign w975[64] = |(datain[55:52] ^ 0);
  assign w975[65] = |(datain[51:48] ^ 0);
  assign w975[66] = |(datain[47:44] ^ 5);
  assign w975[67] = |(datain[43:40] ^ 0);
  assign w975[68] = |(datain[39:36] ^ 12);
  assign w975[69] = |(datain[35:32] ^ 11);
  assign comp[975] = ~(|w975);
  wire [76-1:0] w976;
  assign w976[0] = |(datain[311:308] ^ 13);
  assign w976[1] = |(datain[307:304] ^ 11);
  assign w976[2] = |(datain[303:300] ^ 8);
  assign w976[3] = |(datain[299:296] ^ 14);
  assign w976[4] = |(datain[295:292] ^ 13);
  assign w976[5] = |(datain[291:288] ^ 11);
  assign w976[6] = |(datain[287:284] ^ 8);
  assign w976[7] = |(datain[283:280] ^ 14);
  assign w976[8] = |(datain[279:276] ^ 13);
  assign w976[9] = |(datain[275:272] ^ 3);
  assign w976[10] = |(datain[271:268] ^ 11);
  assign w976[11] = |(datain[267:264] ^ 12);
  assign w976[12] = |(datain[263:260] ^ 0);
  assign w976[13] = |(datain[259:256] ^ 0);
  assign w976[14] = |(datain[255:252] ^ 7);
  assign w976[15] = |(datain[251:248] ^ 12);
  assign w976[16] = |(datain[247:244] ^ 15);
  assign w976[17] = |(datain[243:240] ^ 11);
  assign w976[18] = |(datain[239:236] ^ 10);
  assign w976[19] = |(datain[235:232] ^ 1);
  assign w976[20] = |(datain[231:228] ^ 1);
  assign w976[21] = |(datain[227:224] ^ 3);
  assign w976[22] = |(datain[223:220] ^ 0);
  assign w976[23] = |(datain[219:216] ^ 4);
  assign w976[24] = |(datain[215:212] ^ 2);
  assign w976[25] = |(datain[211:208] ^ 13);
  assign w976[26] = |(datain[207:204] ^ 0);
  assign w976[27] = |(datain[203:200] ^ 5);
  assign w976[28] = |(datain[199:196] ^ 0);
  assign w976[29] = |(datain[195:192] ^ 0);
  assign w976[30] = |(datain[191:188] ^ 10);
  assign w976[31] = |(datain[187:184] ^ 3);
  assign w976[32] = |(datain[183:180] ^ 1);
  assign w976[33] = |(datain[179:176] ^ 3);
  assign w976[34] = |(datain[175:172] ^ 0);
  assign w976[35] = |(datain[171:168] ^ 4);
  assign w976[36] = |(datain[167:164] ^ 11);
  assign w976[37] = |(datain[163:160] ^ 1);
  assign w976[38] = |(datain[159:156] ^ 0);
  assign w976[39] = |(datain[155:152] ^ 6);
  assign w976[40] = |(datain[151:148] ^ 13);
  assign w976[41] = |(datain[147:144] ^ 3);
  assign w976[42] = |(datain[143:140] ^ 14);
  assign w976[43] = |(datain[139:136] ^ 0);
  assign w976[44] = |(datain[135:132] ^ 8);
  assign w976[45] = |(datain[131:128] ^ 14);
  assign w976[46] = |(datain[127:124] ^ 12);
  assign w976[47] = |(datain[123:120] ^ 0);
  assign w976[48] = |(datain[119:116] ^ 11);
  assign w976[49] = |(datain[115:112] ^ 8);
  assign w976[50] = |(datain[111:108] ^ 0);
  assign w976[51] = |(datain[107:104] ^ 9);
  assign w976[52] = |(datain[103:100] ^ 0);
  assign w976[53] = |(datain[99:96] ^ 2);
  assign w976[54] = |(datain[95:92] ^ 11);
  assign w976[55] = |(datain[91:88] ^ 9);
  assign w976[56] = |(datain[87:84] ^ 0);
  assign w976[57] = |(datain[83:80] ^ 2);
  assign w976[58] = |(datain[79:76] ^ 0);
  assign w976[59] = |(datain[75:72] ^ 0);
  assign w976[60] = |(datain[71:68] ^ 11);
  assign w976[61] = |(datain[67:64] ^ 10);
  assign w976[62] = |(datain[63:60] ^ 8);
  assign w976[63] = |(datain[59:56] ^ 0);
  assign w976[64] = |(datain[55:52] ^ 0);
  assign w976[65] = |(datain[51:48] ^ 0);
  assign w976[66] = |(datain[47:44] ^ 12);
  assign w976[67] = |(datain[43:40] ^ 13);
  assign w976[68] = |(datain[39:36] ^ 1);
  assign w976[69] = |(datain[35:32] ^ 3);
  assign w976[70] = |(datain[31:28] ^ 11);
  assign w976[71] = |(datain[27:24] ^ 11);
  assign w976[72] = |(datain[23:20] ^ 7);
  assign w976[73] = |(datain[19:16] ^ 12);
  assign w976[74] = |(datain[15:12] ^ 0);
  assign w976[75] = |(datain[11:8] ^ 1);
  assign comp[976] = ~(|w976);
  wire [44-1:0] w977;
  assign w977[0] = |(datain[311:308] ^ 10);
  assign w977[1] = |(datain[307:304] ^ 1);
  assign w977[2] = |(datain[303:300] ^ 6);
  assign w977[3] = |(datain[299:296] ^ 12);
  assign w977[4] = |(datain[295:292] ^ 0);
  assign w977[5] = |(datain[291:288] ^ 4);
  assign w977[6] = |(datain[287:284] ^ 2);
  assign w977[7] = |(datain[283:280] ^ 6);
  assign w977[8] = |(datain[279:276] ^ 10);
  assign w977[9] = |(datain[275:272] ^ 3);
  assign w977[10] = |(datain[271:268] ^ 12);
  assign w977[11] = |(datain[267:264] ^ 13);
  assign w977[12] = |(datain[263:260] ^ 0);
  assign w977[13] = |(datain[259:256] ^ 4);
  assign w977[14] = |(datain[255:252] ^ 1);
  assign w977[15] = |(datain[251:248] ^ 15);
  assign w977[16] = |(datain[247:244] ^ 0);
  assign w977[17] = |(datain[243:240] ^ 6);
  assign w977[18] = |(datain[239:236] ^ 11);
  assign w977[19] = |(datain[235:232] ^ 8);
  assign w977[20] = |(datain[231:228] ^ 2);
  assign w977[21] = |(datain[227:224] ^ 4);
  assign w977[22] = |(datain[223:220] ^ 3);
  assign w977[23] = |(datain[219:216] ^ 5);
  assign w977[24] = |(datain[215:212] ^ 12);
  assign w977[25] = |(datain[211:208] ^ 13);
  assign w977[26] = |(datain[207:204] ^ 15);
  assign w977[27] = |(datain[203:200] ^ 14);
  assign w977[28] = |(datain[199:196] ^ 8);
  assign w977[29] = |(datain[195:192] ^ 9);
  assign w977[30] = |(datain[191:188] ^ 1);
  assign w977[31] = |(datain[187:184] ^ 14);
  assign w977[32] = |(datain[183:180] ^ 13);
  assign w977[33] = |(datain[179:176] ^ 3);
  assign w977[34] = |(datain[175:172] ^ 0);
  assign w977[35] = |(datain[171:168] ^ 4);
  assign w977[36] = |(datain[167:164] ^ 8);
  assign w977[37] = |(datain[163:160] ^ 12);
  assign w977[38] = |(datain[159:156] ^ 0);
  assign w977[39] = |(datain[155:152] ^ 6);
  assign w977[40] = |(datain[151:148] ^ 13);
  assign w977[41] = |(datain[147:144] ^ 5);
  assign w977[42] = |(datain[143:140] ^ 0);
  assign w977[43] = |(datain[139:136] ^ 4);
  assign comp[977] = ~(|w977);
  wire [28-1:0] w978;
  assign w978[0] = |(datain[311:308] ^ 12);
  assign w978[1] = |(datain[307:304] ^ 13);
  assign w978[2] = |(datain[303:300] ^ 2);
  assign w978[3] = |(datain[299:296] ^ 1);
  assign w978[4] = |(datain[295:292] ^ 8);
  assign w978[5] = |(datain[291:288] ^ 9);
  assign w978[6] = |(datain[287:284] ^ 1);
  assign w978[7] = |(datain[283:280] ^ 14);
  assign w978[8] = |(datain[279:276] ^ 9);
  assign w978[9] = |(datain[275:272] ^ 4);
  assign w978[10] = |(datain[271:268] ^ 0);
  assign w978[11] = |(datain[267:264] ^ 1);
  assign w978[12] = |(datain[263:260] ^ 8);
  assign w978[13] = |(datain[259:256] ^ 12);
  assign w978[14] = |(datain[255:252] ^ 0);
  assign w978[15] = |(datain[251:248] ^ 6);
  assign w978[16] = |(datain[247:244] ^ 9);
  assign w978[17] = |(datain[243:240] ^ 6);
  assign w978[18] = |(datain[239:236] ^ 0);
  assign w978[19] = |(datain[235:232] ^ 1);
  assign w978[20] = |(datain[231:228] ^ 11);
  assign w978[21] = |(datain[227:224] ^ 10);
  assign w978[22] = |(datain[223:220] ^ 8);
  assign w978[23] = |(datain[219:216] ^ 6);
  assign w978[24] = |(datain[215:212] ^ 0);
  assign w978[25] = |(datain[211:208] ^ 1);
  assign w978[26] = |(datain[207:204] ^ 11);
  assign w978[27] = |(datain[203:200] ^ 8);
  assign comp[978] = ~(|w978);
  wire [76-1:0] w979;
  assign w979[0] = |(datain[311:308] ^ 3);
  assign w979[1] = |(datain[307:304] ^ 14);
  assign w979[2] = |(datain[303:300] ^ 8);
  assign w979[3] = |(datain[299:296] ^ 9);
  assign w979[4] = |(datain[295:292] ^ 8);
  assign w979[5] = |(datain[291:288] ^ 6);
  assign w979[6] = |(datain[287:284] ^ 8);
  assign w979[7] = |(datain[283:280] ^ 7);
  assign w979[8] = |(datain[279:276] ^ 0);
  assign w979[9] = |(datain[275:272] ^ 2);
  assign w979[10] = |(datain[271:268] ^ 11);
  assign w979[11] = |(datain[267:264] ^ 8);
  assign w979[12] = |(datain[263:260] ^ 0);
  assign w979[13] = |(datain[259:256] ^ 0);
  assign w979[14] = |(datain[255:252] ^ 4);
  assign w979[15] = |(datain[251:248] ^ 2);
  assign w979[16] = |(datain[247:244] ^ 9);
  assign w979[17] = |(datain[243:240] ^ 9);
  assign w979[18] = |(datain[239:236] ^ 3);
  assign w979[19] = |(datain[235:232] ^ 3);
  assign w979[20] = |(datain[231:228] ^ 12);
  assign w979[21] = |(datain[227:224] ^ 9);
  assign w979[22] = |(datain[223:220] ^ 12);
  assign w979[23] = |(datain[219:216] ^ 13);
  assign w979[24] = |(datain[215:212] ^ 2);
  assign w979[25] = |(datain[211:208] ^ 1);
  assign w979[26] = |(datain[207:204] ^ 11);
  assign w979[27] = |(datain[203:200] ^ 9);
  assign w979[28] = |(datain[199:196] ^ 0);
  assign w979[29] = |(datain[195:192] ^ 3);
  assign w979[30] = |(datain[191:188] ^ 0);
  assign w979[31] = |(datain[187:184] ^ 0);
  assign w979[32] = |(datain[183:180] ^ 11);
  assign w979[33] = |(datain[179:176] ^ 4);
  assign w979[34] = |(datain[175:172] ^ 4);
  assign w979[35] = |(datain[171:168] ^ 0);
  assign w979[36] = |(datain[167:164] ^ 8);
  assign w979[37] = |(datain[163:160] ^ 13);
  assign w979[38] = |(datain[159:156] ^ 9);
  assign w979[39] = |(datain[155:152] ^ 6);
  assign w979[40] = |(datain[151:148] ^ 8);
  assign w979[41] = |(datain[147:144] ^ 6);
  assign w979[42] = |(datain[143:140] ^ 0);
  assign w979[43] = |(datain[139:136] ^ 2);
  assign w979[44] = |(datain[135:132] ^ 12);
  assign w979[45] = |(datain[131:128] ^ 13);
  assign w979[46] = |(datain[127:124] ^ 2);
  assign w979[47] = |(datain[123:120] ^ 1);
  assign w979[48] = |(datain[119:116] ^ 14);
  assign w979[49] = |(datain[115:112] ^ 8);
  assign w979[50] = |(datain[111:108] ^ 6);
  assign w979[51] = |(datain[107:104] ^ 13);
  assign w979[52] = |(datain[103:100] ^ 0);
  assign w979[53] = |(datain[99:96] ^ 0);
  assign w979[54] = |(datain[95:92] ^ 11);
  assign w979[55] = |(datain[91:88] ^ 9);
  assign w979[56] = |(datain[87:84] ^ 9);
  assign w979[57] = |(datain[83:80] ^ 3);
  assign w979[58] = |(datain[79:76] ^ 0);
  assign w979[59] = |(datain[75:72] ^ 1);
  assign w979[60] = |(datain[71:68] ^ 11);
  assign w979[61] = |(datain[67:64] ^ 4);
  assign w979[62] = |(datain[63:60] ^ 4);
  assign w979[63] = |(datain[59:56] ^ 0);
  assign w979[64] = |(datain[55:52] ^ 8);
  assign w979[65] = |(datain[51:48] ^ 13);
  assign w979[66] = |(datain[47:44] ^ 9);
  assign w979[67] = |(datain[43:40] ^ 6);
  assign w979[68] = |(datain[39:36] ^ 0);
  assign w979[69] = |(datain[35:32] ^ 3);
  assign w979[70] = |(datain[31:28] ^ 0);
  assign w979[71] = |(datain[27:24] ^ 1);
  assign w979[72] = |(datain[23:20] ^ 12);
  assign w979[73] = |(datain[19:16] ^ 13);
  assign w979[74] = |(datain[15:12] ^ 2);
  assign w979[75] = |(datain[11:8] ^ 1);
  assign comp[979] = ~(|w979);
  wire [74-1:0] w980;
  assign w980[0] = |(datain[311:308] ^ 8);
  assign w980[1] = |(datain[307:304] ^ 9);
  assign w980[2] = |(datain[303:300] ^ 8);
  assign w980[3] = |(datain[299:296] ^ 6);
  assign w980[4] = |(datain[295:292] ^ 8);
  assign w980[5] = |(datain[291:288] ^ 8);
  assign w980[6] = |(datain[287:284] ^ 0);
  assign w980[7] = |(datain[283:280] ^ 2);
  assign w980[8] = |(datain[279:276] ^ 11);
  assign w980[9] = |(datain[275:272] ^ 8);
  assign w980[10] = |(datain[271:268] ^ 0);
  assign w980[11] = |(datain[267:264] ^ 0);
  assign w980[12] = |(datain[263:260] ^ 4);
  assign w980[13] = |(datain[259:256] ^ 2);
  assign w980[14] = |(datain[255:252] ^ 9);
  assign w980[15] = |(datain[251:248] ^ 9);
  assign w980[16] = |(datain[247:244] ^ 3);
  assign w980[17] = |(datain[243:240] ^ 3);
  assign w980[18] = |(datain[239:236] ^ 12);
  assign w980[19] = |(datain[235:232] ^ 9);
  assign w980[20] = |(datain[231:228] ^ 12);
  assign w980[21] = |(datain[227:224] ^ 13);
  assign w980[22] = |(datain[223:220] ^ 2);
  assign w980[23] = |(datain[219:216] ^ 1);
  assign w980[24] = |(datain[215:212] ^ 11);
  assign w980[25] = |(datain[211:208] ^ 9);
  assign w980[26] = |(datain[207:204] ^ 0);
  assign w980[27] = |(datain[203:200] ^ 3);
  assign w980[28] = |(datain[199:196] ^ 0);
  assign w980[29] = |(datain[195:192] ^ 0);
  assign w980[30] = |(datain[191:188] ^ 11);
  assign w980[31] = |(datain[187:184] ^ 4);
  assign w980[32] = |(datain[183:180] ^ 4);
  assign w980[33] = |(datain[179:176] ^ 0);
  assign w980[34] = |(datain[175:172] ^ 8);
  assign w980[35] = |(datain[171:168] ^ 13);
  assign w980[36] = |(datain[167:164] ^ 9);
  assign w980[37] = |(datain[163:160] ^ 6);
  assign w980[38] = |(datain[159:156] ^ 8);
  assign w980[39] = |(datain[155:152] ^ 7);
  assign w980[40] = |(datain[151:148] ^ 0);
  assign w980[41] = |(datain[147:144] ^ 2);
  assign w980[42] = |(datain[143:140] ^ 12);
  assign w980[43] = |(datain[139:136] ^ 13);
  assign w980[44] = |(datain[135:132] ^ 2);
  assign w980[45] = |(datain[131:128] ^ 1);
  assign w980[46] = |(datain[127:124] ^ 14);
  assign w980[47] = |(datain[123:120] ^ 8);
  assign w980[48] = |(datain[119:116] ^ 6);
  assign w980[49] = |(datain[115:112] ^ 13);
  assign w980[50] = |(datain[111:108] ^ 0);
  assign w980[51] = |(datain[107:104] ^ 0);
  assign w980[52] = |(datain[103:100] ^ 11);
  assign w980[53] = |(datain[99:96] ^ 9);
  assign w980[54] = |(datain[95:92] ^ 9);
  assign w980[55] = |(datain[91:88] ^ 4);
  assign w980[56] = |(datain[87:84] ^ 0);
  assign w980[57] = |(datain[83:80] ^ 1);
  assign w980[58] = |(datain[79:76] ^ 11);
  assign w980[59] = |(datain[75:72] ^ 4);
  assign w980[60] = |(datain[71:68] ^ 4);
  assign w980[61] = |(datain[67:64] ^ 0);
  assign w980[62] = |(datain[63:60] ^ 8);
  assign w980[63] = |(datain[59:56] ^ 13);
  assign w980[64] = |(datain[55:52] ^ 9);
  assign w980[65] = |(datain[51:48] ^ 6);
  assign w980[66] = |(datain[47:44] ^ 0);
  assign w980[67] = |(datain[43:40] ^ 3);
  assign w980[68] = |(datain[39:36] ^ 0);
  assign w980[69] = |(datain[35:32] ^ 1);
  assign w980[70] = |(datain[31:28] ^ 12);
  assign w980[71] = |(datain[27:24] ^ 13);
  assign w980[72] = |(datain[23:20] ^ 2);
  assign w980[73] = |(datain[19:16] ^ 1);
  assign comp[980] = ~(|w980);
  wire [74-1:0] w981;
  assign w981[0] = |(datain[311:308] ^ 0);
  assign w981[1] = |(datain[307:304] ^ 3);
  assign w981[2] = |(datain[303:300] ^ 3);
  assign w981[3] = |(datain[299:296] ^ 2);
  assign w981[4] = |(datain[295:292] ^ 12);
  assign w981[5] = |(datain[291:288] ^ 0);
  assign w981[6] = |(datain[287:284] ^ 14);
  assign w981[7] = |(datain[283:280] ^ 8);
  assign w981[8] = |(datain[279:276] ^ 13);
  assign w981[9] = |(datain[275:272] ^ 13);
  assign w981[10] = |(datain[271:268] ^ 15);
  assign w981[11] = |(datain[267:264] ^ 15);
  assign w981[12] = |(datain[263:260] ^ 11);
  assign w981[13] = |(datain[259:256] ^ 9);
  assign w981[14] = |(datain[255:252] ^ 0);
  assign w981[15] = |(datain[251:248] ^ 3);
  assign w981[16] = |(datain[247:244] ^ 0);
  assign w981[17] = |(datain[243:240] ^ 0);
  assign w981[18] = |(datain[239:236] ^ 11);
  assign w981[19] = |(datain[235:232] ^ 4);
  assign w981[20] = |(datain[231:228] ^ 4);
  assign w981[21] = |(datain[227:224] ^ 0);
  assign w981[22] = |(datain[223:220] ^ 11);
  assign w981[23] = |(datain[219:216] ^ 10);
  assign w981[24] = |(datain[215:212] ^ 2);
  assign w981[25] = |(datain[211:208] ^ 8);
  assign w981[26] = |(datain[207:204] ^ 0);
  assign w981[27] = |(datain[203:200] ^ 3);
  assign w981[28] = |(datain[199:196] ^ 0);
  assign w981[29] = |(datain[195:192] ^ 1);
  assign w981[30] = |(datain[191:188] ^ 14);
  assign w981[31] = |(datain[187:184] ^ 10);
  assign w981[32] = |(datain[183:180] ^ 12);
  assign w981[33] = |(datain[179:176] ^ 13);
  assign w981[34] = |(datain[175:172] ^ 2);
  assign w981[35] = |(datain[171:168] ^ 1);
  assign w981[36] = |(datain[167:164] ^ 11);
  assign w981[37] = |(datain[163:160] ^ 0);
  assign w981[38] = |(datain[159:156] ^ 0);
  assign w981[39] = |(datain[155:152] ^ 2);
  assign w981[40] = |(datain[151:148] ^ 14);
  assign w981[41] = |(datain[147:144] ^ 8);
  assign w981[42] = |(datain[143:140] ^ 12);
  assign w981[43] = |(datain[139:136] ^ 12);
  assign w981[44] = |(datain[135:132] ^ 15);
  assign w981[45] = |(datain[131:128] ^ 15);
  assign w981[46] = |(datain[127:124] ^ 11);
  assign w981[47] = |(datain[123:120] ^ 9);
  assign w981[48] = |(datain[119:116] ^ 2);
  assign w981[49] = |(datain[115:112] ^ 6);
  assign w981[50] = |(datain[111:108] ^ 0);
  assign w981[51] = |(datain[107:104] ^ 2);
  assign w981[52] = |(datain[103:100] ^ 11);
  assign w981[53] = |(datain[99:96] ^ 4);
  assign w981[54] = |(datain[95:92] ^ 4);
  assign w981[55] = |(datain[91:88] ^ 0);
  assign w981[56] = |(datain[87:84] ^ 11);
  assign w981[57] = |(datain[83:80] ^ 10);
  assign w981[58] = |(datain[79:76] ^ 0);
  assign w981[59] = |(datain[75:72] ^ 9);
  assign w981[60] = |(datain[71:68] ^ 0);
  assign w981[61] = |(datain[67:64] ^ 1);
  assign w981[62] = |(datain[63:60] ^ 0);
  assign w981[63] = |(datain[59:56] ^ 1);
  assign w981[64] = |(datain[55:52] ^ 14);
  assign w981[65] = |(datain[51:48] ^ 10);
  assign w981[66] = |(datain[47:44] ^ 12);
  assign w981[67] = |(datain[43:40] ^ 13);
  assign w981[68] = |(datain[39:36] ^ 2);
  assign w981[69] = |(datain[35:32] ^ 1);
  assign w981[70] = |(datain[31:28] ^ 7);
  assign w981[71] = |(datain[27:24] ^ 2);
  assign w981[72] = |(datain[23:20] ^ 10);
  assign w981[73] = |(datain[19:16] ^ 13);
  assign comp[981] = ~(|w981);
  wire [56-1:0] w982;
  assign w982[0] = |(datain[311:308] ^ 12);
  assign w982[1] = |(datain[307:304] ^ 12);
  assign w982[2] = |(datain[303:300] ^ 5);
  assign w982[3] = |(datain[299:296] ^ 13);
  assign w982[4] = |(datain[295:292] ^ 8);
  assign w982[5] = |(datain[291:288] ^ 1);
  assign w982[6] = |(datain[287:284] ^ 14);
  assign w982[7] = |(datain[283:280] ^ 13);
  assign w982[8] = |(datain[279:276] ^ 0);
  assign w982[9] = |(datain[275:272] ^ 6);
  assign w982[10] = |(datain[271:268] ^ 0);
  assign w982[11] = |(datain[267:264] ^ 1);
  assign w982[12] = |(datain[263:260] ^ 12);
  assign w982[13] = |(datain[259:256] ^ 6);
  assign w982[14] = |(datain[255:252] ^ 8);
  assign w982[15] = |(datain[251:248] ^ 6);
  assign w982[16] = |(datain[247:244] ^ 1);
  assign w982[17] = |(datain[243:240] ^ 2);
  assign w982[18] = |(datain[239:236] ^ 0);
  assign w982[19] = |(datain[235:232] ^ 1);
  assign w982[20] = |(datain[231:228] ^ 0);
  assign w982[21] = |(datain[227:224] ^ 1);
  assign w982[22] = |(datain[223:220] ^ 11);
  assign w982[23] = |(datain[219:216] ^ 8);
  assign w982[24] = |(datain[215:212] ^ 0);
  assign w982[25] = |(datain[211:208] ^ 0);
  assign w982[26] = |(datain[207:204] ^ 0);
  assign w982[27] = |(datain[203:200] ^ 0);
  assign w982[28] = |(datain[199:196] ^ 3);
  assign w982[29] = |(datain[195:192] ^ 13);
  assign w982[30] = |(datain[191:188] ^ 0);
  assign w982[31] = |(datain[187:184] ^ 1);
  assign w982[32] = |(datain[183:180] ^ 0);
  assign w982[33] = |(datain[179:176] ^ 0);
  assign w982[34] = |(datain[175:172] ^ 7);
  assign w982[35] = |(datain[171:168] ^ 5);
  assign w982[36] = |(datain[167:164] ^ 0);
  assign w982[37] = |(datain[163:160] ^ 3);
  assign w982[38] = |(datain[159:156] ^ 14);
  assign w982[39] = |(datain[155:152] ^ 9);
  assign w982[40] = |(datain[151:148] ^ 10);
  assign w982[41] = |(datain[147:144] ^ 9);
  assign w982[42] = |(datain[143:140] ^ 0);
  assign w982[43] = |(datain[139:136] ^ 2);
  assign w982[44] = |(datain[135:132] ^ 14);
  assign w982[45] = |(datain[131:128] ^ 8);
  assign w982[46] = |(datain[127:124] ^ 9);
  assign w982[47] = |(datain[123:120] ^ 5);
  assign w982[48] = |(datain[119:116] ^ 0);
  assign w982[49] = |(datain[115:112] ^ 2);
  assign w982[50] = |(datain[111:108] ^ 14);
  assign w982[51] = |(datain[107:104] ^ 8);
  assign w982[52] = |(datain[103:100] ^ 7);
  assign w982[53] = |(datain[99:96] ^ 11);
  assign w982[54] = |(datain[95:92] ^ 0);
  assign w982[55] = |(datain[91:88] ^ 2);
  assign comp[982] = ~(|w982);
  wire [72-1:0] w983;
  assign w983[0] = |(datain[311:308] ^ 8);
  assign w983[1] = |(datain[307:304] ^ 13);
  assign w983[2] = |(datain[303:300] ^ 11);
  assign w983[3] = |(datain[299:296] ^ 6);
  assign w983[4] = |(datain[295:292] ^ 10);
  assign w983[5] = |(datain[291:288] ^ 13);
  assign w983[6] = |(datain[287:284] ^ 0);
  assign w983[7] = |(datain[283:280] ^ 3);
  assign w983[8] = |(datain[279:276] ^ 8);
  assign w983[9] = |(datain[275:272] ^ 11);
  assign w983[10] = |(datain[271:268] ^ 15);
  assign w983[11] = |(datain[267:264] ^ 14);
  assign w983[12] = |(datain[263:260] ^ 10);
  assign w983[13] = |(datain[259:256] ^ 12);
  assign w983[14] = |(datain[255:252] ^ 15);
  assign w983[15] = |(datain[251:248] ^ 6);
  assign w983[16] = |(datain[247:244] ^ 13);
  assign w983[17] = |(datain[243:240] ^ 0);
  assign w983[18] = |(datain[239:236] ^ 10);
  assign w983[19] = |(datain[235:232] ^ 10);
  assign w983[20] = |(datain[231:228] ^ 14);
  assign w983[21] = |(datain[227:224] ^ 2);
  assign w983[22] = |(datain[223:220] ^ 15);
  assign w983[23] = |(datain[219:216] ^ 10);
  assign w983[24] = |(datain[215:212] ^ 12);
  assign w983[25] = |(datain[211:208] ^ 3);
  assign w983[26] = |(datain[207:204] ^ 11);
  assign w983[27] = |(datain[203:200] ^ 4);
  assign w983[28] = |(datain[199:196] ^ 0);
  assign w983[29] = |(datain[195:192] ^ 9);
  assign w983[30] = |(datain[191:188] ^ 8);
  assign w983[31] = |(datain[187:184] ^ 13);
  assign w983[32] = |(datain[183:180] ^ 9);
  assign w983[33] = |(datain[179:176] ^ 6);
  assign w983[34] = |(datain[175:172] ^ 5);
  assign w983[35] = |(datain[171:168] ^ 9);
  assign w983[36] = |(datain[167:164] ^ 0);
  assign w983[37] = |(datain[163:160] ^ 2);
  assign w983[38] = |(datain[159:156] ^ 12);
  assign w983[39] = |(datain[155:152] ^ 13);
  assign w983[40] = |(datain[151:148] ^ 2);
  assign w983[41] = |(datain[147:144] ^ 1);
  assign w983[42] = |(datain[143:140] ^ 15);
  assign w983[43] = |(datain[139:136] ^ 10);
  assign w983[44] = |(datain[135:132] ^ 11);
  assign w983[45] = |(datain[131:128] ^ 8);
  assign w983[46] = |(datain[127:124] ^ 0);
  assign w983[47] = |(datain[123:120] ^ 5);
  assign w983[48] = |(datain[119:116] ^ 2);
  assign w983[49] = |(datain[115:112] ^ 5);
  assign w983[50] = |(datain[111:108] ^ 11);
  assign w983[51] = |(datain[107:104] ^ 11);
  assign w983[52] = |(datain[103:100] ^ 0);
  assign w983[53] = |(datain[99:96] ^ 0);
  assign w983[54] = |(datain[95:92] ^ 11);
  assign w983[55] = |(datain[91:88] ^ 8);
  assign w983[56] = |(datain[87:84] ^ 8);
  assign w983[57] = |(datain[83:80] ^ 14);
  assign w983[58] = |(datain[79:76] ^ 13);
  assign w983[59] = |(datain[75:72] ^ 11);
  assign w983[60] = |(datain[71:68] ^ 11);
  assign w983[61] = |(datain[67:64] ^ 10);
  assign w983[62] = |(datain[63:60] ^ 0);
  assign w983[63] = |(datain[59:56] ^ 0);
  assign w983[64] = |(datain[55:52] ^ 0);
  assign w983[65] = |(datain[51:48] ^ 0);
  assign w983[66] = |(datain[47:44] ^ 12);
  assign w983[67] = |(datain[43:40] ^ 13);
  assign w983[68] = |(datain[39:36] ^ 2);
  assign w983[69] = |(datain[35:32] ^ 1);
  assign w983[70] = |(datain[31:28] ^ 11);
  assign w983[71] = |(datain[27:24] ^ 8);
  assign comp[983] = ~(|w983);
  wire [42-1:0] w984;
  assign w984[0] = |(datain[311:308] ^ 8);
  assign w984[1] = |(datain[307:304] ^ 7);
  assign w984[2] = |(datain[303:300] ^ 0);
  assign w984[3] = |(datain[299:296] ^ 3);
  assign w984[4] = |(datain[295:292] ^ 8);
  assign w984[5] = |(datain[291:288] ^ 13);
  assign w984[6] = |(datain[287:284] ^ 9);
  assign w984[7] = |(datain[283:280] ^ 6);
  assign w984[8] = |(datain[279:276] ^ 0);
  assign w984[9] = |(datain[275:272] ^ 3);
  assign w984[10] = |(datain[271:268] ^ 0);
  assign w984[11] = |(datain[267:264] ^ 1);
  assign w984[12] = |(datain[263:260] ^ 12);
  assign w984[13] = |(datain[259:256] ^ 13);
  assign w984[14] = |(datain[255:252] ^ 2);
  assign w984[15] = |(datain[251:248] ^ 1);
  assign w984[16] = |(datain[247:244] ^ 2);
  assign w984[17] = |(datain[243:240] ^ 14);
  assign w984[18] = |(datain[239:236] ^ 15);
  assign w984[19] = |(datain[235:232] ^ 14);
  assign w984[20] = |(datain[231:228] ^ 0);
  assign w984[21] = |(datain[227:224] ^ 6);
  assign w984[22] = |(datain[223:220] ^ 7);
  assign w984[23] = |(datain[219:216] ^ 2);
  assign w984[24] = |(datain[215:212] ^ 0);
  assign w984[25] = |(datain[211:208] ^ 4);
  assign w984[26] = |(datain[207:204] ^ 14);
  assign w984[27] = |(datain[203:200] ^ 11);
  assign w984[28] = |(datain[199:196] ^ 8);
  assign w984[29] = |(datain[195:192] ^ 9);
  assign w984[30] = |(datain[191:188] ^ 0);
  assign w984[31] = |(datain[187:184] ^ 14);
  assign w984[32] = |(datain[183:180] ^ 14);
  assign w984[33] = |(datain[179:176] ^ 8);
  assign w984[34] = |(datain[175:172] ^ 4);
  assign w984[35] = |(datain[171:168] ^ 9);
  assign w984[36] = |(datain[167:164] ^ 0);
  assign w984[37] = |(datain[163:160] ^ 0);
  assign w984[38] = |(datain[159:156] ^ 11);
  assign w984[39] = |(datain[155:152] ^ 4);
  assign w984[40] = |(datain[151:148] ^ 3);
  assign w984[41] = |(datain[147:144] ^ 11);
  assign comp[984] = ~(|w984);
  wire [30-1:0] w985;
  assign w985[0] = |(datain[311:308] ^ 5);
  assign w985[1] = |(datain[307:304] ^ 10);
  assign w985[2] = |(datain[303:300] ^ 5);
  assign w985[3] = |(datain[299:296] ^ 2);
  assign w985[4] = |(datain[295:292] ^ 8);
  assign w985[5] = |(datain[291:288] ^ 3);
  assign w985[6] = |(datain[287:284] ^ 12);
  assign w985[7] = |(datain[283:280] ^ 2);
  assign w985[8] = |(datain[279:276] ^ 2);
  assign w985[9] = |(datain[275:272] ^ 9);
  assign w985[10] = |(datain[271:268] ^ 11);
  assign w985[11] = |(datain[267:264] ^ 8);
  assign w985[12] = |(datain[263:260] ^ 0);
  assign w985[13] = |(datain[259:256] ^ 2);
  assign w985[14] = |(datain[255:252] ^ 3);
  assign w985[15] = |(datain[251:248] ^ 13);
  assign w985[16] = |(datain[247:244] ^ 12);
  assign w985[17] = |(datain[243:240] ^ 13);
  assign w985[18] = |(datain[239:236] ^ 2);
  assign w985[19] = |(datain[235:232] ^ 1);
  assign w985[20] = |(datain[231:228] ^ 7);
  assign w985[21] = |(datain[227:224] ^ 2);
  assign w985[22] = |(datain[223:220] ^ 7);
  assign w985[23] = |(datain[219:216] ^ 9);
  assign w985[24] = |(datain[215:212] ^ 8);
  assign w985[25] = |(datain[211:208] ^ 11);
  assign w985[26] = |(datain[207:204] ^ 13);
  assign w985[27] = |(datain[203:200] ^ 8);
  assign w985[28] = |(datain[199:196] ^ 5);
  assign w985[29] = |(datain[195:192] ^ 10);
  assign comp[985] = ~(|w985);
  wire [30-1:0] w986;
  assign w986[0] = |(datain[311:308] ^ 0);
  assign w986[1] = |(datain[307:304] ^ 5);
  assign w986[2] = |(datain[303:300] ^ 0);
  assign w986[3] = |(datain[299:296] ^ 3);
  assign w986[4] = |(datain[295:292] ^ 0);
  assign w986[5] = |(datain[291:288] ^ 0);
  assign w986[6] = |(datain[287:284] ^ 5);
  assign w986[7] = |(datain[283:280] ^ 0);
  assign w986[8] = |(datain[279:276] ^ 8);
  assign w986[9] = |(datain[275:272] ^ 11);
  assign w986[10] = |(datain[271:268] ^ 15);
  assign w986[11] = |(datain[267:264] ^ 0);
  assign w986[12] = |(datain[263:260] ^ 11);
  assign w986[13] = |(datain[259:256] ^ 15);
  assign w986[14] = |(datain[255:252] ^ 0);
  assign w986[15] = |(datain[251:248] ^ 0);
  assign w986[16] = |(datain[247:244] ^ 0);
  assign w986[17] = |(datain[243:240] ^ 1);
  assign w986[18] = |(datain[239:236] ^ 11);
  assign w986[19] = |(datain[235:232] ^ 9);
  assign w986[20] = |(datain[231:228] ^ 0);
  assign w986[21] = |(datain[227:224] ^ 5);
  assign w986[22] = |(datain[223:220] ^ 0);
  assign w986[23] = |(datain[219:216] ^ 0);
  assign w986[24] = |(datain[215:212] ^ 15);
  assign w986[25] = |(datain[211:208] ^ 12);
  assign w986[26] = |(datain[207:204] ^ 15);
  assign w986[27] = |(datain[203:200] ^ 3);
  assign w986[28] = |(datain[199:196] ^ 10);
  assign w986[29] = |(datain[195:192] ^ 4);
  assign comp[986] = ~(|w986);
  wire [28-1:0] w987;
  assign w987[0] = |(datain[311:308] ^ 0);
  assign w987[1] = |(datain[307:304] ^ 1);
  assign w987[2] = |(datain[303:300] ^ 10);
  assign w987[3] = |(datain[299:296] ^ 13);
  assign w987[4] = |(datain[295:292] ^ 0);
  assign w987[5] = |(datain[291:288] ^ 5);
  assign w987[6] = |(datain[287:284] ^ 0);
  assign w987[7] = |(datain[283:280] ^ 3);
  assign w987[8] = |(datain[279:276] ^ 0);
  assign w987[9] = |(datain[275:272] ^ 0);
  assign w987[10] = |(datain[271:268] ^ 5);
  assign w987[11] = |(datain[267:264] ^ 0);
  assign w987[12] = |(datain[263:260] ^ 8);
  assign w987[13] = |(datain[259:256] ^ 11);
  assign w987[14] = |(datain[255:252] ^ 15);
  assign w987[15] = |(datain[251:248] ^ 0);
  assign w987[16] = |(datain[247:244] ^ 11);
  assign w987[17] = |(datain[243:240] ^ 15);
  assign w987[18] = |(datain[239:236] ^ 0);
  assign w987[19] = |(datain[235:232] ^ 0);
  assign w987[20] = |(datain[231:228] ^ 0);
  assign w987[21] = |(datain[227:224] ^ 1);
  assign w987[22] = |(datain[223:220] ^ 11);
  assign w987[23] = |(datain[219:216] ^ 9);
  assign w987[24] = |(datain[215:212] ^ 0);
  assign w987[25] = |(datain[211:208] ^ 5);
  assign w987[26] = |(datain[207:204] ^ 0);
  assign w987[27] = |(datain[203:200] ^ 0);
  assign comp[987] = ~(|w987);
  wire [32-1:0] w988;
  assign w988[0] = |(datain[311:308] ^ 12);
  assign w988[1] = |(datain[307:304] ^ 13);
  assign w988[2] = |(datain[303:300] ^ 2);
  assign w988[3] = |(datain[299:296] ^ 1);
  assign w988[4] = |(datain[295:292] ^ 7);
  assign w988[5] = |(datain[291:288] ^ 3);
  assign w988[6] = |(datain[287:284] ^ 0);
  assign w988[7] = |(datain[283:280] ^ 3);
  assign w988[8] = |(datain[279:276] ^ 14);
  assign w988[9] = |(datain[275:272] ^ 9);
  assign w988[10] = |(datain[271:268] ^ 11);
  assign w988[11] = |(datain[267:264] ^ 13);
  assign w988[12] = |(datain[263:260] ^ 0);
  assign w988[13] = |(datain[259:256] ^ 0);
  assign w988[14] = |(datain[255:252] ^ 5);
  assign w988[15] = |(datain[251:248] ^ 14);
  assign w988[16] = |(datain[247:244] ^ 5);
  assign w988[17] = |(datain[243:240] ^ 6);
  assign w988[18] = |(datain[239:236] ^ 8);
  assign w988[19] = |(datain[235:232] ^ 3);
  assign w988[20] = |(datain[231:228] ^ 12);
  assign w988[21] = |(datain[227:224] ^ 6);
  assign w988[22] = |(datain[223:220] ^ 2);
  assign w988[23] = |(datain[219:216] ^ 5);
  assign w988[24] = |(datain[215:212] ^ 10);
  assign w988[25] = |(datain[211:208] ^ 13);
  assign w988[26] = |(datain[207:204] ^ 3);
  assign w988[27] = |(datain[203:200] ^ 13);
  assign w988[28] = |(datain[199:196] ^ 0);
  assign w988[29] = |(datain[195:192] ^ 0);
  assign w988[30] = |(datain[191:188] ^ 15);
  assign w988[31] = |(datain[187:184] ^ 13);
  assign comp[988] = ~(|w988);
  wire [44-1:0] w989;
  assign w989[0] = |(datain[311:308] ^ 0);
  assign w989[1] = |(datain[307:304] ^ 13);
  assign w989[2] = |(datain[303:300] ^ 0);
  assign w989[3] = |(datain[299:296] ^ 0);
  assign w989[4] = |(datain[295:292] ^ 8);
  assign w989[5] = |(datain[291:288] ^ 11);
  assign w989[6] = |(datain[287:284] ^ 15);
  assign w989[7] = |(datain[283:280] ^ 12);
  assign w989[8] = |(datain[279:276] ^ 8);
  assign w989[9] = |(datain[275:272] ^ 13);
  assign w989[10] = |(datain[271:268] ^ 1);
  assign w989[11] = |(datain[267:264] ^ 14);
  assign w989[12] = |(datain[263:260] ^ 2);
  assign w989[13] = |(datain[259:256] ^ 2);
  assign w989[14] = |(datain[255:252] ^ 0);
  assign w989[15] = |(datain[251:248] ^ 0);
  assign w989[16] = |(datain[247:244] ^ 11);
  assign w989[17] = |(datain[243:240] ^ 12);
  assign w989[18] = |(datain[239:236] ^ 4);
  assign w989[19] = |(datain[235:232] ^ 0);
  assign w989[20] = |(datain[231:228] ^ 0);
  assign w989[21] = |(datain[227:224] ^ 0);
  assign w989[22] = |(datain[223:220] ^ 3);
  assign w989[23] = |(datain[219:216] ^ 1);
  assign w989[24] = |(datain[215:212] ^ 2);
  assign w989[25] = |(datain[211:208] ^ 0);
  assign w989[26] = |(datain[207:204] ^ 4);
  assign w989[27] = |(datain[203:200] ^ 3);
  assign w989[28] = |(datain[199:196] ^ 4);
  assign w989[29] = |(datain[195:192] ^ 3);
  assign w989[30] = |(datain[191:188] ^ 4);
  assign w989[31] = |(datain[187:184] ^ 12);
  assign w989[32] = |(datain[183:180] ^ 7);
  assign w989[33] = |(datain[179:176] ^ 5);
  assign w989[34] = |(datain[175:172] ^ 15);
  assign w989[35] = |(datain[171:168] ^ 9);
  assign w989[36] = |(datain[167:164] ^ 12);
  assign w989[37] = |(datain[163:160] ^ 11);
  assign w989[38] = |(datain[159:156] ^ 14);
  assign w989[39] = |(datain[155:152] ^ 7);
  assign w989[40] = |(datain[151:148] ^ 12);
  assign w989[41] = |(datain[147:144] ^ 4);
  assign w989[42] = |(datain[143:140] ^ 0);
  assign w989[43] = |(datain[139:136] ^ 6);
  assign comp[989] = ~(|w989);
  wire [42-1:0] w990;
  assign w990[0] = |(datain[311:308] ^ 7);
  assign w990[1] = |(datain[307:304] ^ 5);
  assign w990[2] = |(datain[303:300] ^ 0);
  assign w990[3] = |(datain[299:296] ^ 3);
  assign w990[4] = |(datain[295:292] ^ 11);
  assign w990[5] = |(datain[291:288] ^ 4);
  assign w990[6] = |(datain[287:284] ^ 15);
  assign w990[7] = |(datain[283:280] ^ 14);
  assign w990[8] = |(datain[279:276] ^ 12);
  assign w990[9] = |(datain[275:272] ^ 15);
  assign w990[10] = |(datain[271:268] ^ 8);
  assign w990[11] = |(datain[267:264] ^ 0);
  assign w990[12] = |(datain[263:260] ^ 15);
  assign w990[13] = |(datain[259:256] ^ 12);
  assign w990[14] = |(datain[255:252] ^ 4);
  assign w990[15] = |(datain[251:248] ^ 11);
  assign w990[16] = |(datain[247:244] ^ 7);
  assign w990[17] = |(datain[243:240] ^ 4);
  assign w990[18] = |(datain[239:236] ^ 0);
  assign w990[19] = |(datain[235:232] ^ 3);
  assign w990[20] = |(datain[231:228] ^ 14);
  assign w990[21] = |(datain[227:224] ^ 9);
  assign w990[22] = |(datain[223:220] ^ 1);
  assign w990[23] = |(datain[219:216] ^ 6);
  assign w990[24] = |(datain[215:212] ^ 0);
  assign w990[25] = |(datain[211:208] ^ 2);
  assign w990[26] = |(datain[207:204] ^ 5);
  assign w990[27] = |(datain[203:200] ^ 0);
  assign w990[28] = |(datain[199:196] ^ 5);
  assign w990[29] = |(datain[195:192] ^ 3);
  assign w990[30] = |(datain[191:188] ^ 5);
  assign w990[31] = |(datain[187:184] ^ 1);
  assign w990[32] = |(datain[183:180] ^ 5);
  assign w990[33] = |(datain[179:176] ^ 2);
  assign w990[34] = |(datain[175:172] ^ 5);
  assign w990[35] = |(datain[171:168] ^ 6);
  assign w990[36] = |(datain[167:164] ^ 5);
  assign w990[37] = |(datain[163:160] ^ 7);
  assign w990[38] = |(datain[159:156] ^ 0);
  assign w990[39] = |(datain[155:152] ^ 6);
  assign w990[40] = |(datain[151:148] ^ 1);
  assign w990[41] = |(datain[147:144] ^ 14);
  assign comp[990] = ~(|w990);
  wire [40-1:0] w991;
  assign w991[0] = |(datain[311:308] ^ 12);
  assign w991[1] = |(datain[307:304] ^ 13);
  assign w991[2] = |(datain[303:300] ^ 2);
  assign w991[3] = |(datain[299:296] ^ 1);
  assign w991[4] = |(datain[295:292] ^ 8);
  assign w991[5] = |(datain[291:288] ^ 1);
  assign w991[6] = |(datain[287:284] ^ 15);
  assign w991[7] = |(datain[283:280] ^ 15);
  assign w991[8] = |(datain[279:276] ^ 12);
  assign w991[9] = |(datain[275:272] ^ 12);
  assign w991[10] = |(datain[271:268] ^ 4);
  assign w991[11] = |(datain[267:264] ^ 4);
  assign w991[12] = |(datain[263:260] ^ 7);
  assign w991[13] = |(datain[259:256] ^ 5);
  assign w991[14] = |(datain[255:252] ^ 0);
  assign w991[15] = |(datain[251:248] ^ 3);
  assign w991[16] = |(datain[247:244] ^ 14);
  assign w991[17] = |(datain[243:240] ^ 9);
  assign w991[18] = |(datain[239:236] ^ 10);
  assign w991[19] = |(datain[235:232] ^ 7);
  assign w991[20] = |(datain[231:228] ^ 0);
  assign w991[21] = |(datain[227:224] ^ 0);
  assign w991[22] = |(datain[223:220] ^ 1);
  assign w991[23] = |(datain[219:216] ^ 14);
  assign w991[24] = |(datain[215:212] ^ 5);
  assign w991[25] = |(datain[211:208] ^ 13);
  assign w991[26] = |(datain[207:204] ^ 4);
  assign w991[27] = |(datain[203:200] ^ 13);
  assign w991[28] = |(datain[199:196] ^ 8);
  assign w991[29] = |(datain[195:192] ^ 14);
  assign w991[30] = |(datain[191:188] ^ 12);
  assign w991[31] = |(datain[187:184] ^ 5);
  assign w991[32] = |(datain[183:180] ^ 8);
  assign w991[33] = |(datain[179:176] ^ 11);
  assign w991[34] = |(datain[175:172] ^ 15);
  assign w991[35] = |(datain[171:168] ^ 3);
  assign w991[36] = |(datain[167:164] ^ 2);
  assign w991[37] = |(datain[163:160] ^ 6);
  assign w991[38] = |(datain[159:156] ^ 8);
  assign w991[39] = |(datain[155:152] ^ 0);
  assign comp[991] = ~(|w991);
  wire [32-1:0] w992;
  assign w992[0] = |(datain[311:308] ^ 4);
  assign w992[1] = |(datain[307:304] ^ 11);
  assign w992[2] = |(datain[303:300] ^ 0);
  assign w992[3] = |(datain[299:296] ^ 0);
  assign w992[4] = |(datain[295:292] ^ 8);
  assign w992[5] = |(datain[291:288] ^ 1);
  assign w992[6] = |(datain[287:284] ^ 12);
  assign w992[7] = |(datain[283:280] ^ 3);
  assign w992[8] = |(datain[279:276] ^ 0);
  assign w992[9] = |(datain[275:272] ^ 0);
  assign w992[10] = |(datain[271:268] ^ 0);
  assign w992[11] = |(datain[267:264] ^ 2);
  assign w992[12] = |(datain[263:260] ^ 14);
  assign w992[13] = |(datain[259:256] ^ 2);
  assign w992[14] = |(datain[255:252] ^ 15);
  assign w992[15] = |(datain[251:248] ^ 4);
  assign w992[16] = |(datain[247:244] ^ 10);
  assign w992[17] = |(datain[243:240] ^ 1);
  assign w992[18] = |(datain[239:236] ^ 1);
  assign w992[19] = |(datain[235:232] ^ 3);
  assign w992[20] = |(datain[231:228] ^ 0);
  assign w992[21] = |(datain[227:224] ^ 4);
  assign w992[22] = |(datain[223:220] ^ 2);
  assign w992[23] = |(datain[219:216] ^ 13);
  assign w992[24] = |(datain[215:212] ^ 0);
  assign w992[25] = |(datain[211:208] ^ 7);
  assign w992[26] = |(datain[207:204] ^ 0);
  assign w992[27] = |(datain[203:200] ^ 0);
  assign w992[28] = |(datain[199:196] ^ 10);
  assign w992[29] = |(datain[195:192] ^ 3);
  assign w992[30] = |(datain[191:188] ^ 1);
  assign w992[31] = |(datain[187:184] ^ 3);
  assign comp[992] = ~(|w992);
  wire [32-1:0] w993;
  assign w993[0] = |(datain[311:308] ^ 15);
  assign w993[1] = |(datain[307:304] ^ 11);
  assign w993[2] = |(datain[303:300] ^ 10);
  assign w993[3] = |(datain[299:296] ^ 0);
  assign w993[4] = |(datain[295:292] ^ 0);
  assign w993[5] = |(datain[291:288] ^ 6);
  assign w993[6] = |(datain[287:284] ^ 7);
  assign w993[7] = |(datain[283:280] ^ 12);
  assign w993[8] = |(datain[279:276] ^ 10);
  assign w993[9] = |(datain[275:272] ^ 2);
  assign w993[10] = |(datain[271:268] ^ 0);
  assign w993[11] = |(datain[267:264] ^ 9);
  assign w993[12] = |(datain[263:260] ^ 7);
  assign w993[13] = |(datain[259:256] ^ 12);
  assign w993[14] = |(datain[255:252] ^ 8);
  assign w993[15] = |(datain[251:248] ^ 11);
  assign w993[16] = |(datain[247:244] ^ 0);
  assign w993[17] = |(datain[243:240] ^ 14);
  assign w993[18] = |(datain[239:236] ^ 0);
  assign w993[19] = |(datain[235:232] ^ 7);
  assign w993[20] = |(datain[231:228] ^ 7);
  assign w993[21] = |(datain[227:224] ^ 12);
  assign w993[22] = |(datain[223:220] ^ 8);
  assign w993[23] = |(datain[219:216] ^ 9);
  assign w993[24] = |(datain[215:212] ^ 0);
  assign w993[25] = |(datain[211:208] ^ 14);
  assign w993[26] = |(datain[207:204] ^ 0);
  assign w993[27] = |(datain[203:200] ^ 10);
  assign w993[28] = |(datain[199:196] ^ 7);
  assign w993[29] = |(datain[195:192] ^ 12);
  assign w993[30] = |(datain[191:188] ^ 14);
  assign w993[31] = |(datain[187:184] ^ 8);
  assign comp[993] = ~(|w993);
  wire [36-1:0] w994;
  assign w994[0] = |(datain[311:308] ^ 10);
  assign w994[1] = |(datain[307:304] ^ 1);
  assign w994[2] = |(datain[303:300] ^ 1);
  assign w994[3] = |(datain[299:296] ^ 3);
  assign w994[4] = |(datain[295:292] ^ 0);
  assign w994[5] = |(datain[291:288] ^ 4);
  assign w994[6] = |(datain[287:284] ^ 2);
  assign w994[7] = |(datain[283:280] ^ 13);
  assign w994[8] = |(datain[279:276] ^ 0);
  assign w994[9] = |(datain[275:272] ^ 7);
  assign w994[10] = |(datain[271:268] ^ 0);
  assign w994[11] = |(datain[267:264] ^ 0);
  assign w994[12] = |(datain[263:260] ^ 10);
  assign w994[13] = |(datain[259:256] ^ 3);
  assign w994[14] = |(datain[255:252] ^ 1);
  assign w994[15] = |(datain[251:248] ^ 3);
  assign w994[16] = |(datain[247:244] ^ 0);
  assign w994[17] = |(datain[243:240] ^ 4);
  assign w994[18] = |(datain[239:236] ^ 11);
  assign w994[19] = |(datain[235:232] ^ 1);
  assign w994[20] = |(datain[231:228] ^ 0);
  assign w994[21] = |(datain[227:224] ^ 6);
  assign w994[22] = |(datain[223:220] ^ 13);
  assign w994[23] = |(datain[219:216] ^ 3);
  assign w994[24] = |(datain[215:212] ^ 14);
  assign w994[25] = |(datain[211:208] ^ 0);
  assign w994[26] = |(datain[207:204] ^ 8);
  assign w994[27] = |(datain[203:200] ^ 14);
  assign w994[28] = |(datain[199:196] ^ 12);
  assign w994[29] = |(datain[195:192] ^ 0);
  assign w994[30] = |(datain[191:188] ^ 11);
  assign w994[31] = |(datain[187:184] ^ 14);
  assign w994[32] = |(datain[183:180] ^ 0);
  assign w994[33] = |(datain[179:176] ^ 0);
  assign w994[34] = |(datain[175:172] ^ 7);
  assign w994[35] = |(datain[171:168] ^ 12);
  assign comp[994] = ~(|w994);
  wire [44-1:0] w995;
  assign w995[0] = |(datain[311:308] ^ 8);
  assign w995[1] = |(datain[307:304] ^ 11);
  assign w995[2] = |(datain[303:300] ^ 14);
  assign w995[3] = |(datain[299:296] ^ 12);
  assign w995[4] = |(datain[295:292] ^ 0);
  assign w995[5] = |(datain[291:288] ^ 14);
  assign w995[6] = |(datain[287:284] ^ 1);
  assign w995[7] = |(datain[283:280] ^ 15);
  assign w995[8] = |(datain[279:276] ^ 11);
  assign w995[9] = |(datain[275:272] ^ 12);
  assign w995[10] = |(datain[271:268] ^ 3);
  assign w995[11] = |(datain[267:264] ^ 4);
  assign w995[12] = |(datain[263:260] ^ 0);
  assign w995[13] = |(datain[259:256] ^ 0);
  assign w995[14] = |(datain[255:252] ^ 15);
  assign w995[15] = |(datain[251:248] ^ 12);
  assign w995[16] = |(datain[247:244] ^ 10);
  assign w995[17] = |(datain[243:240] ^ 13);
  assign w995[18] = |(datain[239:236] ^ 8);
  assign w995[19] = |(datain[235:232] ^ 6);
  assign w995[20] = |(datain[231:228] ^ 12);
  assign w995[21] = |(datain[227:224] ^ 4);
  assign w995[22] = |(datain[223:220] ^ 8);
  assign w995[23] = |(datain[219:216] ^ 9);
  assign w995[24] = |(datain[215:212] ^ 4);
  assign w995[25] = |(datain[211:208] ^ 4);
  assign w995[26] = |(datain[207:204] ^ 15);
  assign w995[27] = |(datain[203:200] ^ 14);
  assign w995[28] = |(datain[199:196] ^ 4);
  assign w995[29] = |(datain[195:192] ^ 4);
  assign w995[30] = |(datain[191:188] ^ 4);
  assign w995[31] = |(datain[187:184] ^ 4);
  assign w995[32] = |(datain[183:180] ^ 8);
  assign w995[33] = |(datain[179:176] ^ 1);
  assign w995[34] = |(datain[175:172] ^ 15);
  assign w995[35] = |(datain[171:168] ^ 12);
  assign w995[36] = |(datain[167:164] ^ 0);
  assign w995[37] = |(datain[163:160] ^ 0);
  assign w995[38] = |(datain[159:156] ^ 0);
  assign w995[39] = |(datain[155:152] ^ 3);
  assign w995[40] = |(datain[151:148] ^ 15);
  assign w995[41] = |(datain[147:144] ^ 2);
  assign w995[42] = |(datain[143:140] ^ 7);
  assign w995[43] = |(datain[139:136] ^ 2);
  assign comp[995] = ~(|w995);
  wire [46-1:0] w996;
  assign w996[0] = |(datain[311:308] ^ 5);
  assign w996[1] = |(datain[307:304] ^ 6);
  assign w996[2] = |(datain[303:300] ^ 5);
  assign w996[3] = |(datain[299:296] ^ 6);
  assign w996[4] = |(datain[295:292] ^ 5);
  assign w996[5] = |(datain[291:288] ^ 6);
  assign w996[6] = |(datain[287:284] ^ 0);
  assign w996[7] = |(datain[283:280] ^ 0);
  assign w996[8] = |(datain[279:276] ^ 0);
  assign w996[9] = |(datain[275:272] ^ 0);
  assign w996[10] = |(datain[271:268] ^ 0);
  assign w996[11] = |(datain[267:264] ^ 0);
  assign w996[12] = |(datain[263:260] ^ 4);
  assign w996[13] = |(datain[259:256] ^ 3);
  assign w996[14] = |(datain[255:252] ^ 4);
  assign w996[15] = |(datain[251:248] ^ 15);
  assign w996[16] = |(datain[247:244] ^ 4);
  assign w996[17] = |(datain[243:240] ^ 13);
  assign w996[18] = |(datain[239:236] ^ 4);
  assign w996[19] = |(datain[235:232] ^ 13);
  assign w996[20] = |(datain[231:228] ^ 4);
  assign w996[21] = |(datain[227:224] ^ 1);
  assign w996[22] = |(datain[223:220] ^ 4);
  assign w996[23] = |(datain[219:216] ^ 14);
  assign w996[24] = |(datain[215:212] ^ 4);
  assign w996[25] = |(datain[211:208] ^ 4);
  assign w996[26] = |(datain[207:204] ^ 2);
  assign w996[27] = |(datain[203:200] ^ 14);
  assign w996[28] = |(datain[199:196] ^ 4);
  assign w996[29] = |(datain[195:192] ^ 3);
  assign w996[30] = |(datain[191:188] ^ 4);
  assign w996[31] = |(datain[187:184] ^ 15);
  assign w996[32] = |(datain[183:180] ^ 4);
  assign w996[33] = |(datain[179:176] ^ 13);
  assign w996[34] = |(datain[175:172] ^ 0);
  assign w996[35] = |(datain[171:168] ^ 0);
  assign w996[36] = |(datain[167:164] ^ 2);
  assign w996[37] = |(datain[163:160] ^ 10);
  assign w996[38] = |(datain[159:156] ^ 2);
  assign w996[39] = |(datain[155:152] ^ 14);
  assign w996[40] = |(datain[151:148] ^ 4);
  assign w996[41] = |(datain[147:144] ^ 3);
  assign w996[42] = |(datain[143:140] ^ 4);
  assign w996[43] = |(datain[139:136] ^ 15);
  assign w996[44] = |(datain[135:132] ^ 4);
  assign w996[45] = |(datain[131:128] ^ 13);
  assign comp[996] = ~(|w996);
  wire [68-1:0] w997;
  assign w997[0] = |(datain[311:308] ^ 0);
  assign w997[1] = |(datain[307:304] ^ 1);
  assign w997[2] = |(datain[303:300] ^ 0);
  assign w997[3] = |(datain[299:296] ^ 2);
  assign w997[4] = |(datain[295:292] ^ 11);
  assign w997[5] = |(datain[291:288] ^ 11);
  assign w997[6] = |(datain[287:284] ^ 0);
  assign w997[7] = |(datain[283:280] ^ 0);
  assign w997[8] = |(datain[279:276] ^ 0);
  assign w997[9] = |(datain[275:272] ^ 2);
  assign w997[10] = |(datain[271:268] ^ 11);
  assign w997[11] = |(datain[267:264] ^ 9);
  assign w997[12] = |(datain[263:260] ^ 0);
  assign w997[13] = |(datain[259:256] ^ 1);
  assign w997[14] = |(datain[255:252] ^ 0);
  assign w997[15] = |(datain[251:248] ^ 0);
  assign w997[16] = |(datain[247:244] ^ 11);
  assign w997[17] = |(datain[243:240] ^ 10);
  assign w997[18] = |(datain[239:236] ^ 8);
  assign w997[19] = |(datain[235:232] ^ 0);
  assign w997[20] = |(datain[231:228] ^ 0);
  assign w997[21] = |(datain[227:224] ^ 0);
  assign w997[22] = |(datain[223:220] ^ 12);
  assign w997[23] = |(datain[219:216] ^ 13);
  assign w997[24] = |(datain[215:212] ^ 1);
  assign w997[25] = |(datain[211:208] ^ 3);
  assign w997[26] = |(datain[207:204] ^ 8);
  assign w997[27] = |(datain[203:200] ^ 1);
  assign w997[28] = |(datain[199:196] ^ 3);
  assign w997[29] = |(datain[195:192] ^ 14);
  assign w997[30] = |(datain[191:188] ^ 10);
  assign w997[31] = |(datain[187:184] ^ 8);
  assign w997[32] = |(datain[183:180] ^ 0);
  assign w997[33] = |(datain[179:176] ^ 3);
  assign w997[34] = |(datain[175:172] ^ 12);
  assign w997[35] = |(datain[171:168] ^ 15);
  assign w997[36] = |(datain[167:164] ^ 12);
  assign w997[37] = |(datain[163:160] ^ 15);
  assign w997[38] = |(datain[159:156] ^ 7);
  assign w997[39] = |(datain[155:152] ^ 4);
  assign w997[40] = |(datain[151:148] ^ 4);
  assign w997[41] = |(datain[147:144] ^ 1);
  assign w997[42] = |(datain[143:140] ^ 11);
  assign w997[43] = |(datain[139:136] ^ 8);
  assign w997[44] = |(datain[135:132] ^ 0);
  assign w997[45] = |(datain[131:128] ^ 1);
  assign w997[46] = |(datain[127:124] ^ 0);
  assign w997[47] = |(datain[123:120] ^ 3);
  assign w997[48] = |(datain[119:116] ^ 11);
  assign w997[49] = |(datain[115:112] ^ 1);
  assign w997[50] = |(datain[111:108] ^ 0);
  assign w997[51] = |(datain[107:104] ^ 3);
  assign w997[52] = |(datain[103:100] ^ 12);
  assign w997[53] = |(datain[99:96] ^ 13);
  assign w997[54] = |(datain[95:92] ^ 1);
  assign w997[55] = |(datain[91:88] ^ 3);
  assign w997[56] = |(datain[87:84] ^ 11);
  assign w997[57] = |(datain[83:80] ^ 15);
  assign w997[58] = |(datain[79:76] ^ 11);
  assign w997[59] = |(datain[75:72] ^ 8);
  assign w997[60] = |(datain[71:68] ^ 0);
  assign w997[61] = |(datain[67:64] ^ 1);
  assign w997[62] = |(datain[63:60] ^ 11);
  assign w997[63] = |(datain[59:56] ^ 14);
  assign w997[64] = |(datain[55:52] ^ 11);
  assign w997[65] = |(datain[51:48] ^ 8);
  assign w997[66] = |(datain[47:44] ^ 0);
  assign w997[67] = |(datain[43:40] ^ 3);
  assign comp[997] = ~(|w997);
  wire [60-1:0] w998;
  assign w998[0] = |(datain[311:308] ^ 0);
  assign w998[1] = |(datain[307:304] ^ 3);
  assign w998[2] = |(datain[303:300] ^ 0);
  assign w998[3] = |(datain[299:296] ^ 0);
  assign w998[4] = |(datain[295:292] ^ 8);
  assign w998[5] = |(datain[291:288] ^ 11);
  assign w998[6] = |(datain[287:284] ^ 15);
  assign w998[7] = |(datain[283:280] ^ 8);
  assign w998[8] = |(datain[279:276] ^ 14);
  assign w998[9] = |(datain[275:272] ^ 11);
  assign w998[10] = |(datain[271:268] ^ 0);
  assign w998[11] = |(datain[267:264] ^ 10);
  assign w998[12] = |(datain[263:260] ^ 3);
  assign w998[13] = |(datain[259:256] ^ 3);
  assign w998[14] = |(datain[255:252] ^ 12);
  assign w998[15] = |(datain[251:248] ^ 0);
  assign w998[16] = |(datain[247:244] ^ 9);
  assign w998[17] = |(datain[243:240] ^ 12);
  assign w998[18] = |(datain[239:236] ^ 2);
  assign w998[19] = |(datain[235:232] ^ 14);
  assign w998[20] = |(datain[231:228] ^ 15);
  assign w998[21] = |(datain[227:224] ^ 15);
  assign w998[22] = |(datain[223:220] ^ 1);
  assign w998[23] = |(datain[219:216] ^ 14);
  assign w998[24] = |(datain[215:212] ^ 0);
  assign w998[25] = |(datain[211:208] ^ 2);
  assign w998[26] = |(datain[207:204] ^ 0);
  assign w998[27] = |(datain[203:200] ^ 2);
  assign w998[28] = |(datain[199:196] ^ 8);
  assign w998[29] = |(datain[195:192] ^ 11);
  assign w998[30] = |(datain[191:188] ^ 12);
  assign w998[31] = |(datain[187:184] ^ 7);
  assign w998[32] = |(datain[183:180] ^ 9);
  assign w998[33] = |(datain[179:176] ^ 12);
  assign w998[34] = |(datain[175:172] ^ 2);
  assign w998[35] = |(datain[171:168] ^ 14);
  assign w998[36] = |(datain[167:164] ^ 15);
  assign w998[37] = |(datain[163:160] ^ 15);
  assign w998[38] = |(datain[159:156] ^ 1);
  assign w998[39] = |(datain[155:152] ^ 14);
  assign w998[40] = |(datain[151:148] ^ 0);
  assign w998[41] = |(datain[147:144] ^ 2);
  assign w998[42] = |(datain[143:140] ^ 0);
  assign w998[43] = |(datain[139:136] ^ 2);
  assign w998[44] = |(datain[135:132] ^ 7);
  assign w998[45] = |(datain[131:128] ^ 3);
  assign w998[46] = |(datain[127:124] ^ 0);
  assign w998[47] = |(datain[123:120] ^ 3);
  assign w998[48] = |(datain[119:116] ^ 4);
  assign w998[49] = |(datain[115:112] ^ 14);
  assign w998[50] = |(datain[111:108] ^ 7);
  assign w998[51] = |(datain[107:104] ^ 5);
  assign w998[52] = |(datain[103:100] ^ 14);
  assign w998[53] = |(datain[99:96] ^ 11);
  assign w998[54] = |(datain[95:92] ^ 8);
  assign w998[55] = |(datain[91:88] ^ 6);
  assign w998[56] = |(datain[87:84] ^ 14);
  assign w998[57] = |(datain[83:80] ^ 14);
  assign w998[58] = |(datain[79:76] ^ 12);
  assign w998[59] = |(datain[75:72] ^ 3);
  assign comp[998] = ~(|w998);
  wire [74-1:0] w999;
  assign w999[0] = |(datain[311:308] ^ 5);
  assign w999[1] = |(datain[307:304] ^ 14);
  assign w999[2] = |(datain[303:300] ^ 8);
  assign w999[3] = |(datain[299:296] ^ 1);
  assign w999[4] = |(datain[295:292] ^ 14);
  assign w999[5] = |(datain[291:288] ^ 14);
  assign w999[6] = |(datain[287:284] ^ 4);
  assign w999[7] = |(datain[283:280] ^ 3);
  assign w999[8] = |(datain[279:276] ^ 0);
  assign w999[9] = |(datain[275:272] ^ 1);
  assign w999[10] = |(datain[271:268] ^ 15);
  assign w999[11] = |(datain[267:264] ^ 10);
  assign w999[12] = |(datain[263:260] ^ 3);
  assign w999[13] = |(datain[259:256] ^ 3);
  assign w999[14] = |(datain[255:252] ^ 12);
  assign w999[15] = |(datain[251:248] ^ 0);
  assign w999[16] = |(datain[247:244] ^ 8);
  assign w999[17] = |(datain[243:240] ^ 14);
  assign w999[18] = |(datain[239:236] ^ 13);
  assign w999[19] = |(datain[235:232] ^ 8);
  assign w999[20] = |(datain[231:228] ^ 8);
  assign w999[21] = |(datain[227:224] ^ 14);
  assign w999[22] = |(datain[223:220] ^ 13);
  assign w999[23] = |(datain[219:216] ^ 0);
  assign w999[24] = |(datain[215:212] ^ 11);
  assign w999[25] = |(datain[211:208] ^ 12);
  assign w999[26] = |(datain[207:204] ^ 0);
  assign w999[27] = |(datain[203:200] ^ 0);
  assign w999[28] = |(datain[199:196] ^ 7);
  assign w999[29] = |(datain[195:192] ^ 12);
  assign w999[30] = |(datain[191:188] ^ 10);
  assign w999[31] = |(datain[187:184] ^ 1);
  assign w999[32] = |(datain[183:180] ^ 1);
  assign w999[33] = |(datain[179:176] ^ 3);
  assign w999[34] = |(datain[175:172] ^ 0);
  assign w999[35] = |(datain[171:168] ^ 4);
  assign w999[36] = |(datain[167:164] ^ 2);
  assign w999[37] = |(datain[163:160] ^ 13);
  assign w999[38] = |(datain[159:156] ^ 0);
  assign w999[39] = |(datain[155:152] ^ 2);
  assign w999[40] = |(datain[151:148] ^ 0);
  assign w999[41] = |(datain[147:144] ^ 0);
  assign w999[42] = |(datain[143:140] ^ 10);
  assign w999[43] = |(datain[139:136] ^ 3);
  assign w999[44] = |(datain[135:132] ^ 1);
  assign w999[45] = |(datain[131:128] ^ 3);
  assign w999[46] = |(datain[127:124] ^ 0);
  assign w999[47] = |(datain[123:120] ^ 4);
  assign w999[48] = |(datain[119:116] ^ 11);
  assign w999[49] = |(datain[115:112] ^ 1);
  assign w999[50] = |(datain[111:108] ^ 0);
  assign w999[51] = |(datain[107:104] ^ 6);
  assign w999[52] = |(datain[103:100] ^ 13);
  assign w999[53] = |(datain[99:96] ^ 3);
  assign w999[54] = |(datain[95:92] ^ 14);
  assign w999[55] = |(datain[91:88] ^ 0);
  assign w999[56] = |(datain[87:84] ^ 8);
  assign w999[57] = |(datain[83:80] ^ 14);
  assign w999[58] = |(datain[79:76] ^ 12);
  assign w999[59] = |(datain[75:72] ^ 0);
  assign w999[60] = |(datain[71:68] ^ 2);
  assign w999[61] = |(datain[67:64] ^ 14);
  assign w999[62] = |(datain[63:60] ^ 8);
  assign w999[63] = |(datain[59:56] ^ 9);
  assign w999[64] = |(datain[55:52] ^ 8);
  assign w999[65] = |(datain[51:48] ^ 4);
  assign w999[66] = |(datain[47:44] ^ 7);
  assign w999[67] = |(datain[43:40] ^ 5);
  assign w999[68] = |(datain[39:36] ^ 0);
  assign w999[69] = |(datain[35:32] ^ 1);
  assign w999[70] = |(datain[31:28] ^ 11);
  assign w999[71] = |(datain[27:24] ^ 15);
  assign w999[72] = |(datain[23:20] ^ 0);
  assign w999[73] = |(datain[19:16] ^ 0);
  assign comp[999] = ~(|w999);
  wire [76-1:0] w1000;
  assign w1000[0] = |(datain[311:308] ^ 1);
  assign w1000[1] = |(datain[307:304] ^ 0);
  assign w1000[2] = |(datain[303:300] ^ 7);
  assign w1000[3] = |(datain[299:296] ^ 5);
  assign w1000[4] = |(datain[295:292] ^ 15);
  assign w1000[5] = |(datain[291:288] ^ 5);
  assign w1000[6] = |(datain[287:284] ^ 3);
  assign w1000[7] = |(datain[283:280] ^ 8);
  assign w1000[8] = |(datain[279:276] ^ 11);
  assign w1000[9] = |(datain[275:272] ^ 15);
  assign w1000[10] = |(datain[271:268] ^ 12);
  assign w1000[11] = |(datain[267:264] ^ 2);
  assign w1000[12] = |(datain[263:260] ^ 0);
  assign w1000[13] = |(datain[259:256] ^ 3);
  assign w1000[14] = |(datain[255:252] ^ 7);
  assign w1000[15] = |(datain[251:248] ^ 5);
  assign w1000[16] = |(datain[247:244] ^ 0);
  assign w1000[17] = |(datain[243:240] ^ 4);
  assign w1000[18] = |(datain[239:236] ^ 8);
  assign w1000[19] = |(datain[235:232] ^ 8);
  assign w1000[20] = |(datain[231:228] ^ 8);
  assign w1000[21] = |(datain[227:224] ^ 15);
  assign w1000[22] = |(datain[223:220] ^ 12);
  assign w1000[23] = |(datain[219:216] ^ 2);
  assign w1000[24] = |(datain[215:212] ^ 0);
  assign w1000[25] = |(datain[211:208] ^ 3);
  assign w1000[26] = |(datain[207:204] ^ 11);
  assign w1000[27] = |(datain[203:200] ^ 3);
  assign w1000[28] = |(datain[199:196] ^ 4);
  assign w1000[29] = |(datain[195:192] ^ 0);
  assign w1000[30] = |(datain[191:188] ^ 8);
  assign w1000[31] = |(datain[187:184] ^ 10);
  assign w1000[32] = |(datain[183:180] ^ 8);
  assign w1000[33] = |(datain[179:176] ^ 7);
  assign w1000[34] = |(datain[175:172] ^ 11);
  assign w1000[35] = |(datain[171:168] ^ 13);
  assign w1000[36] = |(datain[167:164] ^ 0);
  assign w1000[37] = |(datain[163:160] ^ 3);
  assign w1000[38] = |(datain[159:156] ^ 8);
  assign w1000[39] = |(datain[155:152] ^ 8);
  assign w1000[40] = |(datain[151:148] ^ 8);
  assign w1000[41] = |(datain[147:144] ^ 7);
  assign w1000[42] = |(datain[143:140] ^ 11);
  assign w1000[43] = |(datain[139:136] ^ 13);
  assign w1000[44] = |(datain[135:132] ^ 0);
  assign w1000[45] = |(datain[131:128] ^ 1);
  assign w1000[46] = |(datain[127:124] ^ 4);
  assign w1000[47] = |(datain[123:120] ^ 11);
  assign w1000[48] = |(datain[119:116] ^ 7);
  assign w1000[49] = |(datain[115:112] ^ 5);
  assign w1000[50] = |(datain[111:108] ^ 15);
  assign w1000[51] = |(datain[107:104] ^ 5);
  assign w1000[52] = |(datain[103:100] ^ 11);
  assign w1000[53] = |(datain[99:96] ^ 8);
  assign w1000[54] = |(datain[95:92] ^ 0);
  assign w1000[55] = |(datain[91:88] ^ 1);
  assign w1000[56] = |(datain[87:84] ^ 0);
  assign w1000[57] = |(datain[83:80] ^ 3);
  assign w1000[58] = |(datain[79:76] ^ 12);
  assign w1000[59] = |(datain[75:72] ^ 13);
  assign w1000[60] = |(datain[71:68] ^ 1);
  assign w1000[61] = |(datain[67:64] ^ 3);
  assign w1000[62] = |(datain[63:60] ^ 3);
  assign w1000[63] = |(datain[59:56] ^ 1);
  assign w1000[64] = |(datain[55:52] ^ 12);
  assign w1000[65] = |(datain[51:48] ^ 0);
  assign w1000[66] = |(datain[47:44] ^ 8);
  assign w1000[67] = |(datain[43:40] ^ 14);
  assign w1000[68] = |(datain[39:36] ^ 13);
  assign w1000[69] = |(datain[35:32] ^ 8);
  assign w1000[70] = |(datain[31:28] ^ 10);
  assign w1000[71] = |(datain[27:24] ^ 3);
  assign w1000[72] = |(datain[23:20] ^ 8);
  assign w1000[73] = |(datain[19:16] ^ 9);
  assign w1000[74] = |(datain[15:12] ^ 7);
  assign w1000[75] = |(datain[11:8] ^ 12);
  assign comp[1000] = ~(|w1000);
  wire [76-1:0] w1001;
  assign w1001[0] = |(datain[311:308] ^ 7);
  assign w1001[1] = |(datain[307:304] ^ 14);
  assign w1001[2] = |(datain[303:300] ^ 4);
  assign w1001[3] = |(datain[299:296] ^ 1);
  assign w1001[4] = |(datain[295:292] ^ 3);
  assign w1001[5] = |(datain[291:288] ^ 2);
  assign w1001[6] = |(datain[287:284] ^ 15);
  assign w1001[7] = |(datain[283:280] ^ 6);
  assign w1001[8] = |(datain[279:276] ^ 11);
  assign w1001[9] = |(datain[275:272] ^ 2);
  assign w1001[10] = |(datain[271:268] ^ 8);
  assign w1001[11] = |(datain[267:264] ^ 0);
  assign w1001[12] = |(datain[263:260] ^ 12);
  assign w1001[13] = |(datain[259:256] ^ 13);
  assign w1001[14] = |(datain[255:252] ^ 1);
  assign w1001[15] = |(datain[251:248] ^ 3);
  assign w1001[16] = |(datain[247:244] ^ 7);
  assign w1001[17] = |(datain[243:240] ^ 2);
  assign w1001[18] = |(datain[239:236] ^ 14);
  assign w1001[19] = |(datain[235:232] ^ 11);
  assign w1001[20] = |(datain[231:228] ^ 8);
  assign w1001[21] = |(datain[227:224] ^ 0);
  assign w1001[22] = |(datain[223:220] ^ 3);
  assign w1001[23] = |(datain[219:216] ^ 14);
  assign w1001[24] = |(datain[215:212] ^ 2);
  assign w1001[25] = |(datain[211:208] ^ 1);
  assign w1001[26] = |(datain[207:204] ^ 7);
  assign w1001[27] = |(datain[203:200] ^ 14);
  assign w1001[28] = |(datain[199:196] ^ 3);
  assign w1001[29] = |(datain[195:192] ^ 3);
  assign w1001[30] = |(datain[191:188] ^ 7);
  assign w1001[31] = |(datain[187:184] ^ 4);
  assign w1001[32] = |(datain[183:180] ^ 2);
  assign w1001[33] = |(datain[179:176] ^ 8);
  assign w1001[34] = |(datain[175:172] ^ 11);
  assign w1001[35] = |(datain[171:168] ^ 4);
  assign w1001[36] = |(datain[167:164] ^ 0);
  assign w1001[37] = |(datain[163:160] ^ 5);
  assign w1001[38] = |(datain[159:156] ^ 11);
  assign w1001[39] = |(datain[155:152] ^ 1);
  assign w1001[40] = |(datain[151:148] ^ 7);
  assign w1001[41] = |(datain[147:144] ^ 9);
  assign w1001[42] = |(datain[143:140] ^ 12);
  assign w1001[43] = |(datain[139:136] ^ 13);
  assign w1001[44] = |(datain[135:132] ^ 1);
  assign w1001[45] = |(datain[131:128] ^ 6);
  assign w1001[46] = |(datain[127:124] ^ 11);
  assign w1001[47] = |(datain[123:120] ^ 8);
  assign w1001[48] = |(datain[119:116] ^ 0);
  assign w1001[49] = |(datain[115:112] ^ 1);
  assign w1001[50] = |(datain[111:108] ^ 0);
  assign w1001[51] = |(datain[107:104] ^ 3);
  assign w1001[52] = |(datain[103:100] ^ 11);
  assign w1001[53] = |(datain[99:96] ^ 9);
  assign w1001[54] = |(datain[95:92] ^ 0);
  assign w1001[55] = |(datain[91:88] ^ 2);
  assign w1001[56] = |(datain[87:84] ^ 0);
  assign w1001[57] = |(datain[83:80] ^ 0);
  assign w1001[58] = |(datain[79:76] ^ 12);
  assign w1001[59] = |(datain[75:72] ^ 13);
  assign w1001[60] = |(datain[71:68] ^ 1);
  assign w1001[61] = |(datain[67:64] ^ 3);
  assign w1001[62] = |(datain[63:60] ^ 11);
  assign w1001[63] = |(datain[59:56] ^ 4);
  assign w1001[64] = |(datain[55:52] ^ 0);
  assign w1001[65] = |(datain[51:48] ^ 5);
  assign w1001[66] = |(datain[47:44] ^ 11);
  assign w1001[67] = |(datain[43:40] ^ 1);
  assign w1001[68] = |(datain[39:36] ^ 7);
  assign w1001[69] = |(datain[35:32] ^ 9);
  assign w1001[70] = |(datain[31:28] ^ 12);
  assign w1001[71] = |(datain[27:24] ^ 13);
  assign w1001[72] = |(datain[23:20] ^ 1);
  assign w1001[73] = |(datain[19:16] ^ 6);
  assign w1001[74] = |(datain[15:12] ^ 15);
  assign w1001[75] = |(datain[11:8] ^ 12);
  assign comp[1001] = ~(|w1001);
  wire [44-1:0] w1002;
  assign w1002[0] = |(datain[311:308] ^ 0);
  assign w1002[1] = |(datain[307:304] ^ 1);
  assign w1002[2] = |(datain[303:300] ^ 11);
  assign w1002[3] = |(datain[299:296] ^ 14);
  assign w1002[4] = |(datain[295:292] ^ 2);
  assign w1002[5] = |(datain[291:288] ^ 0);
  assign w1002[6] = |(datain[287:284] ^ 7);
  assign w1002[7] = |(datain[283:280] ^ 12);
  assign w1002[8] = |(datain[279:276] ^ 11);
  assign w1002[9] = |(datain[275:272] ^ 9);
  assign w1002[10] = |(datain[271:268] ^ 6);
  assign w1002[11] = |(datain[267:264] ^ 9);
  assign w1002[12] = |(datain[263:260] ^ 0);
  assign w1002[13] = |(datain[259:256] ^ 2);
  assign w1002[14] = |(datain[255:252] ^ 4);
  assign w1002[15] = |(datain[251:248] ^ 1);
  assign w1002[16] = |(datain[247:244] ^ 10);
  assign w1002[17] = |(datain[243:240] ^ 4);
  assign w1002[18] = |(datain[239:236] ^ 14);
  assign w1002[19] = |(datain[235:232] ^ 2);
  assign w1002[20] = |(datain[231:228] ^ 15);
  assign w1002[21] = |(datain[227:224] ^ 13);
  assign w1002[22] = |(datain[223:220] ^ 8);
  assign w1002[23] = |(datain[219:216] ^ 3);
  assign w1002[24] = |(datain[215:212] ^ 2);
  assign w1002[25] = |(datain[211:208] ^ 14);
  assign w1002[26] = |(datain[207:204] ^ 1);
  assign w1002[27] = |(datain[203:200] ^ 3);
  assign w1002[28] = |(datain[199:196] ^ 0);
  assign w1002[29] = |(datain[195:192] ^ 4);
  assign w1002[30] = |(datain[191:188] ^ 1);
  assign w1002[31] = |(datain[187:184] ^ 0);
  assign w1002[32] = |(datain[183:180] ^ 11);
  assign w1002[33] = |(datain[179:176] ^ 11);
  assign w1002[34] = |(datain[175:172] ^ 3);
  assign w1002[35] = |(datain[171:168] ^ 9);
  assign w1002[36] = |(datain[167:164] ^ 0);
  assign w1002[37] = |(datain[163:160] ^ 1);
  assign w1002[38] = |(datain[159:156] ^ 0);
  assign w1002[39] = |(datain[155:152] ^ 6);
  assign w1002[40] = |(datain[151:148] ^ 5);
  assign w1002[41] = |(datain[147:144] ^ 3);
  assign w1002[42] = |(datain[143:140] ^ 12);
  assign w1002[43] = |(datain[139:136] ^ 11);
  assign comp[1002] = ~(|w1002);
  wire [46-1:0] w1003;
  assign w1003[0] = |(datain[311:308] ^ 0);
  assign w1003[1] = |(datain[307:304] ^ 1);
  assign w1003[2] = |(datain[303:300] ^ 8);
  assign w1003[3] = |(datain[299:296] ^ 11);
  assign w1003[4] = |(datain[295:292] ^ 15);
  assign w1003[5] = |(datain[291:288] ^ 14);
  assign w1003[6] = |(datain[287:284] ^ 8);
  assign w1003[7] = |(datain[283:280] ^ 13);
  assign w1003[8] = |(datain[279:276] ^ 1);
  assign w1003[9] = |(datain[275:272] ^ 6);
  assign w1003[10] = |(datain[271:268] ^ 1);
  assign w1003[11] = |(datain[267:264] ^ 15);
  assign w1003[12] = |(datain[263:260] ^ 0);
  assign w1003[13] = |(datain[259:256] ^ 1);
  assign w1003[14] = |(datain[255:252] ^ 8);
  assign w1003[15] = |(datain[251:248] ^ 13);
  assign w1003[16] = |(datain[247:244] ^ 0);
  assign w1003[17] = |(datain[243:240] ^ 14);
  assign w1003[18] = |(datain[239:236] ^ 2);
  assign w1003[19] = |(datain[235:232] ^ 15);
  assign w1003[20] = |(datain[231:228] ^ 0);
  assign w1003[21] = |(datain[227:224] ^ 14);
  assign w1003[22] = |(datain[223:220] ^ 2);
  assign w1003[23] = |(datain[219:216] ^ 11);
  assign w1003[24] = |(datain[215:212] ^ 12);
  assign w1003[25] = |(datain[211:208] ^ 10);
  assign w1003[26] = |(datain[207:204] ^ 15);
  assign w1003[27] = |(datain[203:200] ^ 12);
  assign w1003[28] = |(datain[199:196] ^ 10);
  assign w1003[29] = |(datain[195:192] ^ 12);
  assign w1003[30] = |(datain[191:188] ^ 13);
  assign w1003[31] = |(datain[187:184] ^ 0);
  assign w1003[32] = |(datain[183:180] ^ 12);
  assign w1003[33] = |(datain[179:176] ^ 8);
  assign w1003[34] = |(datain[175:172] ^ 10);
  assign w1003[35] = |(datain[171:168] ^ 10);
  assign w1003[36] = |(datain[167:164] ^ 14);
  assign w1003[37] = |(datain[163:160] ^ 2);
  assign w1003[38] = |(datain[159:156] ^ 15);
  assign w1003[39] = |(datain[155:152] ^ 10);
  assign w1003[40] = |(datain[151:148] ^ 14);
  assign w1003[41] = |(datain[147:144] ^ 9);
  assign w1003[42] = |(datain[143:140] ^ 4);
  assign w1003[43] = |(datain[139:136] ^ 8);
  assign w1003[44] = |(datain[135:132] ^ 0);
  assign w1003[45] = |(datain[131:128] ^ 12);
  assign comp[1003] = ~(|w1003);
  wire [42-1:0] w1004;
  assign w1004[0] = |(datain[311:308] ^ 0);
  assign w1004[1] = |(datain[307:304] ^ 1);
  assign w1004[2] = |(datain[303:300] ^ 8);
  assign w1004[3] = |(datain[299:296] ^ 11);
  assign w1004[4] = |(datain[295:292] ^ 15);
  assign w1004[5] = |(datain[291:288] ^ 14);
  assign w1004[6] = |(datain[287:284] ^ 8);
  assign w1004[7] = |(datain[283:280] ^ 13);
  assign w1004[8] = |(datain[279:276] ^ 1);
  assign w1004[9] = |(datain[275:272] ^ 6);
  assign w1004[10] = |(datain[271:268] ^ 1);
  assign w1004[11] = |(datain[267:264] ^ 15);
  assign w1004[12] = |(datain[263:260] ^ 0);
  assign w1004[13] = |(datain[259:256] ^ 1);
  assign w1004[14] = |(datain[255:252] ^ 8);
  assign w1004[15] = |(datain[251:248] ^ 13);
  assign w1004[16] = |(datain[247:244] ^ 0);
  assign w1004[17] = |(datain[243:240] ^ 14);
  assign w1004[18] = |(datain[239:236] ^ 2);
  assign w1004[19] = |(datain[235:232] ^ 15);
  assign w1004[20] = |(datain[231:228] ^ 0);
  assign w1004[21] = |(datain[227:224] ^ 14);
  assign w1004[22] = |(datain[223:220] ^ 2);
  assign w1004[23] = |(datain[219:216] ^ 11);
  assign w1004[24] = |(datain[215:212] ^ 12);
  assign w1004[25] = |(datain[211:208] ^ 10);
  assign w1004[26] = |(datain[207:204] ^ 15);
  assign w1004[27] = |(datain[203:200] ^ 12);
  assign w1004[28] = |(datain[199:196] ^ 10);
  assign w1004[29] = |(datain[195:192] ^ 12);
  assign w1004[30] = |(datain[191:188] ^ 13);
  assign w1004[31] = |(datain[187:184] ^ 0);
  assign w1004[32] = |(datain[183:180] ^ 12);
  assign w1004[33] = |(datain[179:176] ^ 8);
  assign w1004[34] = |(datain[175:172] ^ 10);
  assign w1004[35] = |(datain[171:168] ^ 10);
  assign w1004[36] = |(datain[167:164] ^ 14);
  assign w1004[37] = |(datain[163:160] ^ 2);
  assign w1004[38] = |(datain[159:156] ^ 15);
  assign w1004[39] = |(datain[155:152] ^ 10);
  assign w1004[40] = |(datain[151:148] ^ 14);
  assign w1004[41] = |(datain[147:144] ^ 9);
  assign comp[1004] = ~(|w1004);
  wire [42-1:0] w1005;
  assign w1005[0] = |(datain[311:308] ^ 1);
  assign w1005[1] = |(datain[307:304] ^ 10);
  assign w1005[2] = |(datain[303:300] ^ 7);
  assign w1005[3] = |(datain[299:296] ^ 2);
  assign w1005[4] = |(datain[295:292] ^ 2);
  assign w1005[5] = |(datain[291:288] ^ 1);
  assign w1005[6] = |(datain[287:284] ^ 8);
  assign w1005[7] = |(datain[283:280] ^ 0);
  assign w1005[8] = |(datain[279:276] ^ 15);
  assign w1005[9] = |(datain[275:272] ^ 14);
  assign w1005[10] = |(datain[271:268] ^ 0);
  assign w1005[11] = |(datain[267:264] ^ 2);
  assign w1005[12] = |(datain[263:260] ^ 7);
  assign w1005[13] = |(datain[259:256] ^ 5);
  assign w1005[14] = |(datain[255:252] ^ 1);
  assign w1005[15] = |(datain[251:248] ^ 12);
  assign w1005[16] = |(datain[247:244] ^ 11);
  assign w1005[17] = |(datain[243:240] ^ 4);
  assign w1005[18] = |(datain[239:236] ^ 2);
  assign w1005[19] = |(datain[235:232] ^ 12);
  assign w1005[20] = |(datain[231:228] ^ 12);
  assign w1005[21] = |(datain[227:224] ^ 13);
  assign w1005[22] = |(datain[223:220] ^ 2);
  assign w1005[23] = |(datain[219:216] ^ 1);
  assign w1005[24] = |(datain[215:212] ^ 8);
  assign w1005[25] = |(datain[211:208] ^ 3);
  assign w1005[26] = |(datain[207:204] ^ 15);
  assign w1005[27] = |(datain[203:200] ^ 10);
  assign w1005[28] = |(datain[199:196] ^ 3);
  assign w1005[29] = |(datain[195:192] ^ 12);
  assign w1005[30] = |(datain[191:188] ^ 7);
  assign w1005[31] = |(datain[187:184] ^ 15);
  assign w1005[32] = |(datain[183:180] ^ 1);
  assign w1005[33] = |(datain[179:176] ^ 3);
  assign w1005[34] = |(datain[175:172] ^ 8);
  assign w1005[35] = |(datain[171:168] ^ 13);
  assign w1005[36] = |(datain[167:164] ^ 7);
  assign w1005[37] = |(datain[163:160] ^ 6);
  assign w1005[38] = |(datain[159:156] ^ 0);
  assign w1005[39] = |(datain[155:152] ^ 7);
  assign w1005[40] = |(datain[151:148] ^ 15);
  assign w1005[41] = |(datain[147:144] ^ 12);
  assign comp[1005] = ~(|w1005);
  wire [24-1:0] w1006;
  assign w1006[0] = |(datain[311:308] ^ 11);
  assign w1006[1] = |(datain[307:304] ^ 4);
  assign w1006[2] = |(datain[303:300] ^ 4);
  assign w1006[3] = |(datain[299:296] ^ 14);
  assign w1006[4] = |(datain[295:292] ^ 12);
  assign w1006[5] = |(datain[291:288] ^ 13);
  assign w1006[6] = |(datain[287:284] ^ 2);
  assign w1006[7] = |(datain[283:280] ^ 1);
  assign w1006[8] = |(datain[279:276] ^ 7);
  assign w1006[9] = |(datain[275:272] ^ 2);
  assign w1006[10] = |(datain[271:268] ^ 0);
  assign w1006[11] = |(datain[267:264] ^ 15);
  assign w1006[12] = |(datain[263:260] ^ 11);
  assign w1006[13] = |(datain[259:256] ^ 10);
  assign w1006[14] = |(datain[255:252] ^ 9);
  assign w1006[15] = |(datain[251:248] ^ 14);
  assign w1006[16] = |(datain[247:244] ^ 0);
  assign w1006[17] = |(datain[243:240] ^ 0);
  assign w1006[18] = |(datain[239:236] ^ 11);
  assign w1006[19] = |(datain[235:232] ^ 8);
  assign w1006[20] = |(datain[231:228] ^ 0);
  assign w1006[21] = |(datain[227:224] ^ 2);
  assign w1006[22] = |(datain[223:220] ^ 3);
  assign w1006[23] = |(datain[219:216] ^ 13);
  assign comp[1006] = ~(|w1006);
  wire [44-1:0] w1007;
  assign w1007[0] = |(datain[311:308] ^ 1);
  assign w1007[1] = |(datain[307:304] ^ 14);
  assign w1007[2] = |(datain[303:300] ^ 7);
  assign w1007[3] = |(datain[299:296] ^ 12);
  assign w1007[4] = |(datain[295:292] ^ 0);
  assign w1007[5] = |(datain[291:288] ^ 15);
  assign w1007[6] = |(datain[287:284] ^ 11);
  assign w1007[7] = |(datain[283:280] ^ 4);
  assign w1007[8] = |(datain[279:276] ^ 1);
  assign w1007[9] = |(datain[275:272] ^ 3);
  assign w1007[10] = |(datain[271:268] ^ 12);
  assign w1007[11] = |(datain[267:264] ^ 13);
  assign w1007[12] = |(datain[263:260] ^ 2);
  assign w1007[13] = |(datain[259:256] ^ 15);
  assign w1007[14] = |(datain[255:252] ^ 1);
  assign w1007[15] = |(datain[251:248] ^ 14);
  assign w1007[16] = |(datain[247:244] ^ 5);
  assign w1007[17] = |(datain[243:240] ^ 2);
  assign w1007[18] = |(datain[239:236] ^ 11);
  assign w1007[19] = |(datain[235:232] ^ 4);
  assign w1007[20] = |(datain[231:228] ^ 1);
  assign w1007[21] = |(datain[227:224] ^ 3);
  assign w1007[22] = |(datain[223:220] ^ 12);
  assign w1007[23] = |(datain[219:216] ^ 13);
  assign w1007[24] = |(datain[215:212] ^ 2);
  assign w1007[25] = |(datain[211:208] ^ 15);
  assign w1007[26] = |(datain[207:204] ^ 5);
  assign w1007[27] = |(datain[203:200] ^ 10);
  assign w1007[28] = |(datain[199:196] ^ 0);
  assign w1007[29] = |(datain[195:192] ^ 7);
  assign w1007[30] = |(datain[191:188] ^ 14);
  assign w1007[31] = |(datain[187:184] ^ 11);
  assign w1007[32] = |(datain[183:180] ^ 0);
  assign w1007[33] = |(datain[179:176] ^ 5);
  assign w1007[34] = |(datain[175:172] ^ 9);
  assign w1007[35] = |(datain[171:168] ^ 0);
  assign w1007[36] = |(datain[167:164] ^ 12);
  assign w1007[37] = |(datain[163:160] ^ 4);
  assign w1007[38] = |(datain[159:156] ^ 1);
  assign w1007[39] = |(datain[155:152] ^ 6);
  assign w1007[40] = |(datain[151:148] ^ 4);
  assign w1007[41] = |(datain[147:144] ^ 12);
  assign w1007[42] = |(datain[143:140] ^ 0);
  assign w1007[43] = |(datain[139:136] ^ 0);
  assign comp[1007] = ~(|w1007);
  wire [32-1:0] w1008;
  assign w1008[0] = |(datain[311:308] ^ 14);
  assign w1008[1] = |(datain[307:304] ^ 2);
  assign w1008[2] = |(datain[303:300] ^ 15);
  assign w1008[3] = |(datain[299:296] ^ 10);
  assign w1008[4] = |(datain[295:292] ^ 8);
  assign w1008[5] = |(datain[291:288] ^ 11);
  assign w1008[6] = |(datain[287:284] ^ 13);
  assign w1008[7] = |(datain[283:280] ^ 7);
  assign w1008[8] = |(datain[279:276] ^ 12);
  assign w1008[9] = |(datain[275:272] ^ 3);
  assign w1008[10] = |(datain[271:268] ^ 11);
  assign w1008[11] = |(datain[267:264] ^ 4);
  assign w1008[12] = |(datain[263:260] ^ 4);
  assign w1008[13] = |(datain[259:256] ^ 0);
  assign w1008[14] = |(datain[255:252] ^ 11);
  assign w1008[15] = |(datain[251:248] ^ 9);
  assign w1008[16] = |(datain[247:244] ^ 15);
  assign w1008[17] = |(datain[243:240] ^ 13);
  assign w1008[18] = |(datain[239:236] ^ 0);
  assign w1008[19] = |(datain[235:232] ^ 7);
  assign w1008[20] = |(datain[231:228] ^ 11);
  assign w1008[21] = |(datain[227:224] ^ 10);
  assign w1008[22] = |(datain[223:220] ^ 0);
  assign w1008[23] = |(datain[219:216] ^ 0);
  assign w1008[24] = |(datain[215:212] ^ 0);
  assign w1008[25] = |(datain[211:208] ^ 1);
  assign w1008[26] = |(datain[207:204] ^ 14);
  assign w1008[27] = |(datain[203:200] ^ 11);
  assign w1008[28] = |(datain[199:196] ^ 4);
  assign w1008[29] = |(datain[195:192] ^ 15);
  assign w1008[30] = |(datain[191:188] ^ 11);
  assign w1008[31] = |(datain[187:184] ^ 8);
  assign comp[1008] = ~(|w1008);
  wire [20-1:0] w1009;
  assign w1009[0] = |(datain[311:308] ^ 4);
  assign w1009[1] = |(datain[307:304] ^ 11);
  assign w1009[2] = |(datain[303:300] ^ 12);
  assign w1009[3] = |(datain[299:296] ^ 13);
  assign w1009[4] = |(datain[295:292] ^ 2);
  assign w1009[5] = |(datain[291:288] ^ 1);
  assign w1009[6] = |(datain[287:284] ^ 7);
  assign w1009[7] = |(datain[283:280] ^ 2);
  assign w1009[8] = |(datain[279:276] ^ 0);
  assign w1009[9] = |(datain[275:272] ^ 3);
  assign w1009[10] = |(datain[271:268] ^ 14);
  assign w1009[11] = |(datain[267:264] ^ 9);
  assign w1009[12] = |(datain[263:260] ^ 13);
  assign w1009[13] = |(datain[259:256] ^ 7);
  assign w1009[14] = |(datain[255:252] ^ 0);
  assign w1009[15] = |(datain[251:248] ^ 0);
  assign w1009[16] = |(datain[247:244] ^ 5);
  assign w1009[17] = |(datain[243:240] ^ 14);
  assign w1009[18] = |(datain[239:236] ^ 5);
  assign w1009[19] = |(datain[235:232] ^ 6);
  assign comp[1009] = ~(|w1009);
  wire [74-1:0] w1010;
  assign w1010[0] = |(datain[311:308] ^ 8);
  assign w1010[1] = |(datain[307:304] ^ 9);
  assign w1010[2] = |(datain[303:300] ^ 1);
  assign w1010[3] = |(datain[299:296] ^ 6);
  assign w1010[4] = |(datain[295:292] ^ 14);
  assign w1010[5] = |(datain[291:288] ^ 5);
  assign w1010[6] = |(datain[287:284] ^ 0);
  assign w1010[7] = |(datain[283:280] ^ 3);
  assign w1010[8] = |(datain[279:276] ^ 11);
  assign w1010[9] = |(datain[275:272] ^ 0);
  assign w1010[10] = |(datain[271:268] ^ 0);
  assign w1010[11] = |(datain[267:264] ^ 0);
  assign w1010[12] = |(datain[263:260] ^ 14);
  assign w1010[13] = |(datain[259:256] ^ 8);
  assign w1010[14] = |(datain[255:252] ^ 14);
  assign w1010[15] = |(datain[251:248] ^ 11);
  assign w1010[16] = |(datain[247:244] ^ 15);
  assign w1010[17] = |(datain[243:240] ^ 14);
  assign w1010[18] = |(datain[239:236] ^ 11);
  assign w1010[19] = |(datain[235:232] ^ 4);
  assign w1010[20] = |(datain[231:228] ^ 4);
  assign w1010[21] = |(datain[227:224] ^ 0);
  assign w1010[22] = |(datain[223:220] ^ 11);
  assign w1010[23] = |(datain[219:216] ^ 9);
  assign w1010[24] = |(datain[215:212] ^ 1);
  assign w1010[25] = |(datain[211:208] ^ 8);
  assign w1010[26] = |(datain[207:204] ^ 0);
  assign w1010[27] = |(datain[203:200] ^ 0);
  assign w1010[28] = |(datain[199:196] ^ 11);
  assign w1010[29] = |(datain[195:192] ^ 10);
  assign w1010[30] = |(datain[191:188] ^ 14);
  assign w1010[31] = |(datain[187:184] ^ 3);
  assign w1010[32] = |(datain[183:180] ^ 0);
  assign w1010[33] = |(datain[179:176] ^ 3);
  assign w1010[34] = |(datain[175:172] ^ 12);
  assign w1010[35] = |(datain[171:168] ^ 13);
  assign w1010[36] = |(datain[167:164] ^ 5);
  assign w1010[37] = |(datain[163:160] ^ 0);
  assign w1010[38] = |(datain[159:156] ^ 11);
  assign w1010[39] = |(datain[155:152] ^ 0);
  assign w1010[40] = |(datain[151:148] ^ 0);
  assign w1010[41] = |(datain[147:144] ^ 2);
  assign w1010[42] = |(datain[143:140] ^ 14);
  assign w1010[43] = |(datain[139:136] ^ 8);
  assign w1010[44] = |(datain[135:132] ^ 13);
  assign w1010[45] = |(datain[131:128] ^ 12);
  assign w1010[46] = |(datain[127:124] ^ 15);
  assign w1010[47] = |(datain[123:120] ^ 14);
  assign w1010[48] = |(datain[119:116] ^ 0);
  assign w1010[49] = |(datain[115:112] ^ 14);
  assign w1010[50] = |(datain[111:108] ^ 1);
  assign w1010[51] = |(datain[107:104] ^ 15);
  assign w1010[52] = |(datain[103:100] ^ 11);
  assign w1010[53] = |(datain[99:96] ^ 4);
  assign w1010[54] = |(datain[95:92] ^ 4);
  assign w1010[55] = |(datain[91:88] ^ 0);
  assign w1010[56] = |(datain[87:84] ^ 11);
  assign w1010[57] = |(datain[83:80] ^ 9);
  assign w1010[58] = |(datain[79:76] ^ 15);
  assign w1010[59] = |(datain[75:72] ^ 15);
  assign w1010[60] = |(datain[71:68] ^ 0);
  assign w1010[61] = |(datain[67:64] ^ 1);
  assign w1010[62] = |(datain[63:60] ^ 11);
  assign w1010[63] = |(datain[59:56] ^ 10);
  assign w1010[64] = |(datain[55:52] ^ 0);
  assign w1010[65] = |(datain[51:48] ^ 0);
  assign w1010[66] = |(datain[47:44] ^ 0);
  assign w1010[67] = |(datain[43:40] ^ 2);
  assign w1010[68] = |(datain[39:36] ^ 12);
  assign w1010[69] = |(datain[35:32] ^ 13);
  assign w1010[70] = |(datain[31:28] ^ 5);
  assign w1010[71] = |(datain[27:24] ^ 0);
  assign w1010[72] = |(datain[23:20] ^ 5);
  assign w1010[73] = |(datain[19:16] ^ 10);
  assign comp[1010] = ~(|w1010);
  wire [74-1:0] w1011;
  assign w1011[0] = |(datain[311:308] ^ 8);
  assign w1011[1] = |(datain[307:304] ^ 9);
  assign w1011[2] = |(datain[303:300] ^ 1);
  assign w1011[3] = |(datain[299:296] ^ 6);
  assign w1011[4] = |(datain[295:292] ^ 14);
  assign w1011[5] = |(datain[291:288] ^ 5);
  assign w1011[6] = |(datain[287:284] ^ 0);
  assign w1011[7] = |(datain[283:280] ^ 3);
  assign w1011[8] = |(datain[279:276] ^ 11);
  assign w1011[9] = |(datain[275:272] ^ 0);
  assign w1011[10] = |(datain[271:268] ^ 0);
  assign w1011[11] = |(datain[267:264] ^ 0);
  assign w1011[12] = |(datain[263:260] ^ 14);
  assign w1011[13] = |(datain[259:256] ^ 8);
  assign w1011[14] = |(datain[255:252] ^ 0);
  assign w1011[15] = |(datain[251:248] ^ 5);
  assign w1011[16] = |(datain[247:244] ^ 15);
  assign w1011[17] = |(datain[243:240] ^ 15);
  assign w1011[18] = |(datain[239:236] ^ 11);
  assign w1011[19] = |(datain[235:232] ^ 4);
  assign w1011[20] = |(datain[231:228] ^ 4);
  assign w1011[21] = |(datain[227:224] ^ 0);
  assign w1011[22] = |(datain[223:220] ^ 11);
  assign w1011[23] = |(datain[219:216] ^ 9);
  assign w1011[24] = |(datain[215:212] ^ 1);
  assign w1011[25] = |(datain[211:208] ^ 8);
  assign w1011[26] = |(datain[207:204] ^ 0);
  assign w1011[27] = |(datain[203:200] ^ 0);
  assign w1011[28] = |(datain[199:196] ^ 11);
  assign w1011[29] = |(datain[195:192] ^ 10);
  assign w1011[30] = |(datain[191:188] ^ 14);
  assign w1011[31] = |(datain[187:184] ^ 3);
  assign w1011[32] = |(datain[183:180] ^ 0);
  assign w1011[33] = |(datain[179:176] ^ 3);
  assign w1011[34] = |(datain[175:172] ^ 12);
  assign w1011[35] = |(datain[171:168] ^ 13);
  assign w1011[36] = |(datain[167:164] ^ 5);
  assign w1011[37] = |(datain[163:160] ^ 0);
  assign w1011[38] = |(datain[159:156] ^ 11);
  assign w1011[39] = |(datain[155:152] ^ 0);
  assign w1011[40] = |(datain[151:148] ^ 0);
  assign w1011[41] = |(datain[147:144] ^ 2);
  assign w1011[42] = |(datain[143:140] ^ 14);
  assign w1011[43] = |(datain[139:136] ^ 8);
  assign w1011[44] = |(datain[135:132] ^ 15);
  assign w1011[45] = |(datain[131:128] ^ 6);
  assign w1011[46] = |(datain[127:124] ^ 15);
  assign w1011[47] = |(datain[123:120] ^ 14);
  assign w1011[48] = |(datain[119:116] ^ 0);
  assign w1011[49] = |(datain[115:112] ^ 14);
  assign w1011[50] = |(datain[111:108] ^ 1);
  assign w1011[51] = |(datain[107:104] ^ 15);
  assign w1011[52] = |(datain[103:100] ^ 11);
  assign w1011[53] = |(datain[99:96] ^ 4);
  assign w1011[54] = |(datain[95:92] ^ 4);
  assign w1011[55] = |(datain[91:88] ^ 0);
  assign w1011[56] = |(datain[87:84] ^ 11);
  assign w1011[57] = |(datain[83:80] ^ 9);
  assign w1011[58] = |(datain[79:76] ^ 2);
  assign w1011[59] = |(datain[75:72] ^ 11);
  assign w1011[60] = |(datain[71:68] ^ 0);
  assign w1011[61] = |(datain[67:64] ^ 2);
  assign w1011[62] = |(datain[63:60] ^ 11);
  assign w1011[63] = |(datain[59:56] ^ 10);
  assign w1011[64] = |(datain[55:52] ^ 0);
  assign w1011[65] = |(datain[51:48] ^ 0);
  assign w1011[66] = |(datain[47:44] ^ 0);
  assign w1011[67] = |(datain[43:40] ^ 2);
  assign w1011[68] = |(datain[39:36] ^ 12);
  assign w1011[69] = |(datain[35:32] ^ 13);
  assign w1011[70] = |(datain[31:28] ^ 5);
  assign w1011[71] = |(datain[27:24] ^ 0);
  assign w1011[72] = |(datain[23:20] ^ 5);
  assign w1011[73] = |(datain[19:16] ^ 10);
  assign comp[1011] = ~(|w1011);
  wire [64-1:0] w1012;
  assign w1012[0] = |(datain[311:308] ^ 11);
  assign w1012[1] = |(datain[307:304] ^ 4);
  assign w1012[2] = |(datain[303:300] ^ 1);
  assign w1012[3] = |(datain[299:296] ^ 10);
  assign w1012[4] = |(datain[295:292] ^ 12);
  assign w1012[5] = |(datain[291:288] ^ 13);
  assign w1012[6] = |(datain[287:284] ^ 2);
  assign w1012[7] = |(datain[283:280] ^ 1);
  assign w1012[8] = |(datain[279:276] ^ 8);
  assign w1012[9] = |(datain[275:272] ^ 11);
  assign w1012[10] = |(datain[271:268] ^ 2);
  assign w1012[11] = |(datain[267:264] ^ 14);
  assign w1012[12] = |(datain[263:260] ^ 2);
  assign w1012[13] = |(datain[259:256] ^ 12);
  assign w1012[14] = |(datain[255:252] ^ 0);
  assign w1012[15] = |(datain[251:248] ^ 1);
  assign w1012[16] = |(datain[247:244] ^ 11);
  assign w1012[17] = |(datain[243:240] ^ 10);
  assign w1012[18] = |(datain[239:236] ^ 14);
  assign w1012[19] = |(datain[235:232] ^ 6);
  assign w1012[20] = |(datain[231:228] ^ 0);
  assign w1012[21] = |(datain[227:224] ^ 2);
  assign w1012[22] = |(datain[223:220] ^ 11);
  assign w1012[23] = |(datain[219:216] ^ 8);
  assign w1012[24] = |(datain[215:212] ^ 2);
  assign w1012[25] = |(datain[211:208] ^ 4);
  assign w1012[26] = |(datain[207:204] ^ 2);
  assign w1012[27] = |(datain[203:200] ^ 5);
  assign w1012[28] = |(datain[199:196] ^ 12);
  assign w1012[29] = |(datain[195:192] ^ 13);
  assign w1012[30] = |(datain[191:188] ^ 2);
  assign w1012[31] = |(datain[187:184] ^ 1);
  assign w1012[32] = |(datain[183:180] ^ 11);
  assign w1012[33] = |(datain[179:176] ^ 4);
  assign w1012[34] = |(datain[175:172] ^ 2);
  assign w1012[35] = |(datain[171:168] ^ 10);
  assign w1012[36] = |(datain[167:164] ^ 12);
  assign w1012[37] = |(datain[163:160] ^ 13);
  assign w1012[38] = |(datain[159:156] ^ 2);
  assign w1012[39] = |(datain[155:152] ^ 1);
  assign w1012[40] = |(datain[151:148] ^ 8);
  assign w1012[41] = |(datain[147:144] ^ 0);
  assign w1012[42] = |(datain[143:140] ^ 15);
  assign w1012[43] = |(datain[139:136] ^ 10);
  assign w1012[44] = |(datain[135:132] ^ 0);
  assign w1012[45] = |(datain[131:128] ^ 11);
  assign w1012[46] = |(datain[127:124] ^ 7);
  assign w1012[47] = |(datain[123:120] ^ 4);
  assign w1012[48] = |(datain[119:116] ^ 0);
  assign w1012[49] = |(datain[115:112] ^ 7);
  assign w1012[50] = |(datain[111:108] ^ 8);
  assign w1012[51] = |(datain[107:104] ^ 0);
  assign w1012[52] = |(datain[103:100] ^ 15);
  assign w1012[53] = |(datain[99:96] ^ 10);
  assign w1012[54] = |(datain[95:92] ^ 1);
  assign w1012[55] = |(datain[91:88] ^ 7);
  assign w1012[56] = |(datain[87:84] ^ 7);
  assign w1012[57] = |(datain[83:80] ^ 4);
  assign w1012[58] = |(datain[79:76] ^ 0);
  assign w1012[59] = |(datain[75:72] ^ 2);
  assign w1012[60] = |(datain[71:68] ^ 14);
  assign w1012[61] = |(datain[67:64] ^ 11);
  assign w1012[62] = |(datain[63:60] ^ 0);
  assign w1012[63] = |(datain[59:56] ^ 11);
  assign comp[1012] = ~(|w1012);
  wire [42-1:0] w1013;
  assign w1013[0] = |(datain[311:308] ^ 14);
  assign w1013[1] = |(datain[307:304] ^ 12);
  assign w1013[2] = |(datain[303:300] ^ 0);
  assign w1013[3] = |(datain[299:296] ^ 1);
  assign w1013[4] = |(datain[295:292] ^ 11);
  assign w1013[5] = |(datain[291:288] ^ 10);
  assign w1013[6] = |(datain[287:284] ^ 1);
  assign w1013[7] = |(datain[283:280] ^ 4);
  assign w1013[8] = |(datain[279:276] ^ 15);
  assign w1013[9] = |(datain[275:272] ^ 13);
  assign w1013[10] = |(datain[271:268] ^ 12);
  assign w1013[11] = |(datain[267:264] ^ 13);
  assign w1013[12] = |(datain[263:260] ^ 2);
  assign w1013[13] = |(datain[259:256] ^ 1);
  assign w1013[14] = |(datain[255:252] ^ 7);
  assign w1013[15] = |(datain[251:248] ^ 2);
  assign w1013[16] = |(datain[247:244] ^ 1);
  assign w1013[17] = |(datain[243:240] ^ 3);
  assign w1013[18] = |(datain[239:236] ^ 3);
  assign w1013[19] = |(datain[235:232] ^ 3);
  assign w1013[20] = |(datain[231:228] ^ 13);
  assign w1013[21] = |(datain[227:224] ^ 2);
  assign w1013[22] = |(datain[223:220] ^ 3);
  assign w1013[23] = |(datain[219:216] ^ 3);
  assign w1013[24] = |(datain[215:212] ^ 12);
  assign w1013[25] = |(datain[211:208] ^ 9);
  assign w1013[26] = |(datain[207:204] ^ 11);
  assign w1013[27] = |(datain[203:200] ^ 8);
  assign w1013[28] = |(datain[199:196] ^ 0);
  assign w1013[29] = |(datain[195:192] ^ 0);
  assign w1013[30] = |(datain[191:188] ^ 4);
  assign w1013[31] = |(datain[187:184] ^ 2);
  assign w1013[32] = |(datain[183:180] ^ 12);
  assign w1013[33] = |(datain[179:176] ^ 13);
  assign w1013[34] = |(datain[175:172] ^ 2);
  assign w1013[35] = |(datain[171:168] ^ 1);
  assign w1013[36] = |(datain[167:164] ^ 11);
  assign w1013[37] = |(datain[163:160] ^ 4);
  assign w1013[38] = |(datain[159:156] ^ 4);
  assign w1013[39] = |(datain[155:152] ^ 0);
  assign w1013[40] = |(datain[151:148] ^ 11);
  assign w1013[41] = |(datain[147:144] ^ 10);
  assign comp[1013] = ~(|w1013);
  wire [30-1:0] w1014;
  assign w1014[0] = |(datain[311:308] ^ 15);
  assign w1014[1] = |(datain[307:304] ^ 15);
  assign w1014[2] = |(datain[303:300] ^ 14);
  assign w1014[3] = |(datain[299:296] ^ 8);
  assign w1014[4] = |(datain[295:292] ^ 14);
  assign w1014[5] = |(datain[291:288] ^ 7);
  assign w1014[6] = |(datain[287:284] ^ 15);
  assign w1014[7] = |(datain[283:280] ^ 15);
  assign w1014[8] = |(datain[279:276] ^ 7);
  assign w1014[9] = |(datain[275:272] ^ 4);
  assign w1014[10] = |(datain[271:268] ^ 2);
  assign w1014[11] = |(datain[267:264] ^ 5);
  assign w1014[12] = |(datain[263:260] ^ 2);
  assign w1014[13] = |(datain[259:256] ^ 14);
  assign w1014[14] = |(datain[255:252] ^ 12);
  assign w1014[15] = |(datain[251:248] ^ 6);
  assign w1014[16] = |(datain[247:244] ^ 0);
  assign w1014[17] = |(datain[243:240] ^ 6);
  assign w1014[18] = |(datain[239:236] ^ 2);
  assign w1014[19] = |(datain[235:232] ^ 9);
  assign w1014[20] = |(datain[231:228] ^ 0);
  assign w1014[21] = |(datain[227:224] ^ 1);
  assign w1014[22] = |(datain[223:220] ^ 0);
  assign w1014[23] = |(datain[219:216] ^ 0);
  assign w1014[24] = |(datain[215:212] ^ 11);
  assign w1014[25] = |(datain[211:208] ^ 8);
  assign w1014[26] = |(datain[207:204] ^ 0);
  assign w1014[27] = |(datain[203:200] ^ 1);
  assign w1014[28] = |(datain[199:196] ^ 0);
  assign w1014[29] = |(datain[195:192] ^ 3);
  assign comp[1014] = ~(|w1014);
  wire [46-1:0] w1015;
  assign w1015[0] = |(datain[311:308] ^ 12);
  assign w1015[1] = |(datain[307:304] ^ 13);
  assign w1015[2] = |(datain[303:300] ^ 2);
  assign w1015[3] = |(datain[299:296] ^ 1);
  assign w1015[4] = |(datain[295:292] ^ 11);
  assign w1015[5] = |(datain[291:288] ^ 9);
  assign w1015[6] = |(datain[287:284] ^ 0);
  assign w1015[7] = |(datain[283:280] ^ 7);
  assign w1015[8] = |(datain[279:276] ^ 0);
  assign w1015[9] = |(datain[275:272] ^ 0);
  assign w1015[10] = |(datain[271:268] ^ 11);
  assign w1015[11] = |(datain[267:264] ^ 15);
  assign w1015[12] = |(datain[263:260] ^ 0);
  assign w1015[13] = |(datain[259:256] ^ 3);
  assign w1015[14] = |(datain[255:252] ^ 0);
  assign w1015[15] = |(datain[251:248] ^ 1);
  assign w1015[16] = |(datain[247:244] ^ 8);
  assign w1015[17] = |(datain[243:240] ^ 11);
  assign w1015[18] = |(datain[239:236] ^ 3);
  assign w1015[19] = |(datain[235:232] ^ 5);
  assign w1015[20] = |(datain[231:228] ^ 8);
  assign w1015[21] = |(datain[227:224] ^ 1);
  assign w1015[22] = |(datain[223:220] ^ 12);
  assign w1015[23] = |(datain[219:216] ^ 6);
  assign w1015[24] = |(datain[215:212] ^ 9);
  assign w1015[25] = |(datain[211:208] ^ 10);
  assign w1015[26] = |(datain[207:204] ^ 0);
  assign w1015[27] = |(datain[203:200] ^ 3);
  assign w1015[28] = |(datain[199:196] ^ 11);
  assign w1015[29] = |(datain[195:192] ^ 15);
  assign w1015[30] = |(datain[191:188] ^ 0);
  assign w1015[31] = |(datain[187:184] ^ 0);
  assign w1015[32] = |(datain[183:180] ^ 0);
  assign w1015[33] = |(datain[179:176] ^ 1);
  assign w1015[34] = |(datain[175:172] ^ 15);
  assign w1015[35] = |(datain[171:168] ^ 12);
  assign w1015[36] = |(datain[167:164] ^ 15);
  assign w1015[37] = |(datain[163:160] ^ 3);
  assign w1015[38] = |(datain[159:156] ^ 10);
  assign w1015[39] = |(datain[155:152] ^ 4);
  assign w1015[40] = |(datain[151:148] ^ 14);
  assign w1015[41] = |(datain[147:144] ^ 11);
  assign w1015[42] = |(datain[143:140] ^ 2);
  assign w1015[43] = |(datain[139:136] ^ 2);
  assign w1015[44] = |(datain[135:132] ^ 9);
  assign w1015[45] = |(datain[131:128] ^ 0);
  assign comp[1015] = ~(|w1015);
  wire [74-1:0] w1016;
  assign w1016[0] = |(datain[311:308] ^ 0);
  assign w1016[1] = |(datain[307:304] ^ 1);
  assign w1016[2] = |(datain[303:300] ^ 0);
  assign w1016[3] = |(datain[299:296] ^ 3);
  assign w1016[4] = |(datain[295:292] ^ 11);
  assign w1016[5] = |(datain[291:288] ^ 10);
  assign w1016[6] = |(datain[287:284] ^ 0);
  assign w1016[7] = |(datain[283:280] ^ 0);
  assign w1016[8] = |(datain[279:276] ^ 0);
  assign w1016[9] = |(datain[275:272] ^ 0);
  assign w1016[10] = |(datain[271:268] ^ 11);
  assign w1016[11] = |(datain[267:264] ^ 9);
  assign w1016[12] = |(datain[263:260] ^ 0);
  assign w1016[13] = |(datain[259:256] ^ 1);
  assign w1016[14] = |(datain[255:252] ^ 0);
  assign w1016[15] = |(datain[251:248] ^ 0);
  assign w1016[16] = |(datain[247:244] ^ 11);
  assign w1016[17] = |(datain[243:240] ^ 11);
  assign w1016[18] = |(datain[239:236] ^ 10);
  assign w1016[19] = |(datain[235:232] ^ 0);
  assign w1016[20] = |(datain[231:228] ^ 0);
  assign w1016[21] = |(datain[227:224] ^ 1);
  assign w1016[22] = |(datain[223:220] ^ 12);
  assign w1016[23] = |(datain[219:216] ^ 13);
  assign w1016[24] = |(datain[215:212] ^ 1);
  assign w1016[25] = |(datain[211:208] ^ 3);
  assign w1016[26] = |(datain[207:204] ^ 7);
  assign w1016[27] = |(datain[203:200] ^ 2);
  assign w1016[28] = |(datain[199:196] ^ 1);
  assign w1016[29] = |(datain[195:192] ^ 5);
  assign w1016[30] = |(datain[191:188] ^ 11);
  assign w1016[31] = |(datain[187:184] ^ 8);
  assign w1016[32] = |(datain[183:180] ^ 0);
  assign w1016[33] = |(datain[179:176] ^ 2);
  assign w1016[34] = |(datain[175:172] ^ 0);
  assign w1016[35] = |(datain[171:168] ^ 3);
  assign w1016[36] = |(datain[167:164] ^ 11);
  assign w1016[37] = |(datain[163:160] ^ 10);
  assign w1016[38] = |(datain[159:156] ^ 0);
  assign w1016[39] = |(datain[155:152] ^ 0);
  assign w1016[40] = |(datain[151:148] ^ 0);
  assign w1016[41] = |(datain[147:144] ^ 0);
  assign w1016[42] = |(datain[143:140] ^ 11);
  assign w1016[43] = |(datain[139:136] ^ 9);
  assign w1016[44] = |(datain[135:132] ^ 0);
  assign w1016[45] = |(datain[131:128] ^ 8);
  assign w1016[46] = |(datain[127:124] ^ 0);
  assign w1016[47] = |(datain[123:120] ^ 0);
  assign w1016[48] = |(datain[119:116] ^ 11);
  assign w1016[49] = |(datain[115:112] ^ 11);
  assign w1016[50] = |(datain[111:108] ^ 10);
  assign w1016[51] = |(datain[107:104] ^ 0);
  assign w1016[52] = |(datain[103:100] ^ 0);
  assign w1016[53] = |(datain[99:96] ^ 3);
  assign w1016[54] = |(datain[95:92] ^ 12);
  assign w1016[55] = |(datain[91:88] ^ 13);
  assign w1016[56] = |(datain[87:84] ^ 1);
  assign w1016[57] = |(datain[83:80] ^ 3);
  assign w1016[58] = |(datain[79:76] ^ 7);
  assign w1016[59] = |(datain[75:72] ^ 2);
  assign w1016[60] = |(datain[71:68] ^ 0);
  assign w1016[61] = |(datain[67:64] ^ 5);
  assign w1016[62] = |(datain[63:60] ^ 11);
  assign w1016[63] = |(datain[59:56] ^ 8);
  assign w1016[64] = |(datain[55:52] ^ 0);
  assign w1016[65] = |(datain[51:48] ^ 0);
  assign w1016[66] = |(datain[47:44] ^ 4);
  assign w1016[67] = |(datain[43:40] ^ 12);
  assign w1016[68] = |(datain[39:36] ^ 12);
  assign w1016[69] = |(datain[35:32] ^ 13);
  assign w1016[70] = |(datain[31:28] ^ 2);
  assign w1016[71] = |(datain[27:24] ^ 1);
  assign w1016[72] = |(datain[23:20] ^ 0);
  assign w1016[73] = |(datain[19:16] ^ 14);
  assign comp[1016] = ~(|w1016);
  wire [74-1:0] w1017;
  assign w1017[0] = |(datain[311:308] ^ 8);
  assign w1017[1] = |(datain[307:304] ^ 11);
  assign w1017[2] = |(datain[303:300] ^ 12);
  assign w1017[3] = |(datain[299:296] ^ 10);
  assign w1017[4] = |(datain[295:292] ^ 11);
  assign w1017[5] = |(datain[291:288] ^ 4);
  assign w1017[6] = |(datain[287:284] ^ 3);
  assign w1017[7] = |(datain[283:280] ^ 15);
  assign w1017[8] = |(datain[279:276] ^ 12);
  assign w1017[9] = |(datain[275:272] ^ 13);
  assign w1017[10] = |(datain[271:268] ^ 2);
  assign w1017[11] = |(datain[267:264] ^ 1);
  assign w1017[12] = |(datain[263:260] ^ 5);
  assign w1017[13] = |(datain[259:256] ^ 0);
  assign w1017[14] = |(datain[255:252] ^ 5);
  assign w1017[15] = |(datain[251:248] ^ 2);
  assign w1017[16] = |(datain[247:244] ^ 14);
  assign w1017[17] = |(datain[243:240] ^ 8);
  assign w1017[18] = |(datain[239:236] ^ 11);
  assign w1017[19] = |(datain[235:232] ^ 14);
  assign w1017[20] = |(datain[231:228] ^ 0);
  assign w1017[21] = |(datain[227:224] ^ 1);
  assign w1017[22] = |(datain[223:220] ^ 5);
  assign w1017[23] = |(datain[219:216] ^ 10);
  assign w1017[24] = |(datain[215:212] ^ 5);
  assign w1017[25] = |(datain[211:208] ^ 9);
  assign w1017[26] = |(datain[207:204] ^ 11);
  assign w1017[27] = |(datain[203:200] ^ 4);
  assign w1017[28] = |(datain[199:196] ^ 4);
  assign w1017[29] = |(datain[195:192] ^ 0);
  assign w1017[30] = |(datain[191:188] ^ 12);
  assign w1017[31] = |(datain[187:184] ^ 13);
  assign w1017[32] = |(datain[183:180] ^ 2);
  assign w1017[33] = |(datain[179:176] ^ 1);
  assign w1017[34] = |(datain[175:172] ^ 5);
  assign w1017[35] = |(datain[171:168] ^ 10);
  assign w1017[36] = |(datain[167:164] ^ 7);
  assign w1017[37] = |(datain[163:160] ^ 2);
  assign w1017[38] = |(datain[159:156] ^ 1);
  assign w1017[39] = |(datain[155:152] ^ 11);
  assign w1017[40] = |(datain[151:148] ^ 3);
  assign w1017[41] = |(datain[147:144] ^ 3);
  assign w1017[42] = |(datain[143:140] ^ 12);
  assign w1017[43] = |(datain[139:136] ^ 9);
  assign w1017[44] = |(datain[135:132] ^ 11);
  assign w1017[45] = |(datain[131:128] ^ 8);
  assign w1017[46] = |(datain[127:124] ^ 0);
  assign w1017[47] = |(datain[123:120] ^ 0);
  assign w1017[48] = |(datain[119:116] ^ 4);
  assign w1017[49] = |(datain[115:112] ^ 2);
  assign w1017[50] = |(datain[111:108] ^ 12);
  assign w1017[51] = |(datain[107:104] ^ 13);
  assign w1017[52] = |(datain[103:100] ^ 2);
  assign w1017[53] = |(datain[99:96] ^ 1);
  assign w1017[54] = |(datain[95:92] ^ 11);
  assign w1017[55] = |(datain[91:88] ^ 4);
  assign w1017[56] = |(datain[87:84] ^ 4);
  assign w1017[57] = |(datain[83:80] ^ 0);
  assign w1017[58] = |(datain[79:76] ^ 12);
  assign w1017[59] = |(datain[75:72] ^ 13);
  assign w1017[60] = |(datain[71:68] ^ 2);
  assign w1017[61] = |(datain[67:64] ^ 1);
  assign w1017[62] = |(datain[63:60] ^ 8);
  assign w1017[63] = |(datain[59:56] ^ 11);
  assign w1017[64] = |(datain[55:52] ^ 12);
  assign w1017[65] = |(datain[51:48] ^ 14);
  assign w1017[66] = |(datain[47:44] ^ 8);
  assign w1017[67] = |(datain[43:40] ^ 11);
  assign w1017[68] = |(datain[39:36] ^ 13);
  assign w1017[69] = |(datain[35:32] ^ 7);
  assign w1017[70] = |(datain[31:28] ^ 8);
  assign w1017[71] = |(datain[27:24] ^ 0);
  assign w1017[72] = |(datain[23:20] ^ 15);
  assign w1017[73] = |(datain[19:16] ^ 1);
  assign comp[1017] = ~(|w1017);
  wire [74-1:0] w1018;
  assign w1018[0] = |(datain[311:308] ^ 0);
  assign w1018[1] = |(datain[307:304] ^ 6);
  assign w1018[2] = |(datain[303:300] ^ 11);
  assign w1018[3] = |(datain[299:296] ^ 7);
  assign w1018[4] = |(datain[295:292] ^ 0);
  assign w1018[5] = |(datain[291:288] ^ 3);
  assign w1018[6] = |(datain[287:284] ^ 14);
  assign w1018[7] = |(datain[283:280] ^ 9);
  assign w1018[8] = |(datain[279:276] ^ 10);
  assign w1018[9] = |(datain[275:272] ^ 3);
  assign w1018[10] = |(datain[271:268] ^ 11);
  assign w1018[11] = |(datain[267:264] ^ 8);
  assign w1018[12] = |(datain[263:260] ^ 0);
  assign w1018[13] = |(datain[259:256] ^ 3);
  assign w1018[14] = |(datain[255:252] ^ 11);
  assign w1018[15] = |(datain[251:248] ^ 4);
  assign w1018[16] = |(datain[247:244] ^ 4);
  assign w1018[17] = |(datain[243:240] ^ 0);
  assign w1018[18] = |(datain[239:236] ^ 11);
  assign w1018[19] = |(datain[235:232] ^ 9);
  assign w1018[20] = |(datain[231:228] ^ 13);
  assign w1018[21] = |(datain[227:224] ^ 7);
  assign w1018[22] = |(datain[223:220] ^ 0);
  assign w1018[23] = |(datain[219:216] ^ 1);
  assign w1018[24] = |(datain[215:212] ^ 11);
  assign w1018[25] = |(datain[211:208] ^ 10);
  assign w1018[26] = |(datain[207:204] ^ 14);
  assign w1018[27] = |(datain[203:200] ^ 0);
  assign w1018[28] = |(datain[199:196] ^ 0);
  assign w1018[29] = |(datain[195:192] ^ 1);
  assign w1018[30] = |(datain[191:188] ^ 12);
  assign w1018[31] = |(datain[187:184] ^ 13);
  assign w1018[32] = |(datain[183:180] ^ 2);
  assign w1018[33] = |(datain[179:176] ^ 1);
  assign w1018[34] = |(datain[175:172] ^ 3);
  assign w1018[35] = |(datain[171:168] ^ 3);
  assign w1018[36] = |(datain[167:164] ^ 14);
  assign w1018[37] = |(datain[163:160] ^ 13);
  assign w1018[38] = |(datain[159:156] ^ 2);
  assign w1018[39] = |(datain[155:152] ^ 6);
  assign w1018[40] = |(datain[151:148] ^ 8);
  assign w1018[41] = |(datain[147:144] ^ 9);
  assign w1018[42] = |(datain[143:140] ^ 6);
  assign w1018[43] = |(datain[139:136] ^ 13);
  assign w1018[44] = |(datain[135:132] ^ 1);
  assign w1018[45] = |(datain[131:128] ^ 5);
  assign w1018[46] = |(datain[127:124] ^ 2);
  assign w1018[47] = |(datain[123:120] ^ 6);
  assign w1018[48] = |(datain[119:116] ^ 8);
  assign w1018[49] = |(datain[115:112] ^ 9);
  assign w1018[50] = |(datain[111:108] ^ 6);
  assign w1018[51] = |(datain[107:104] ^ 13);
  assign w1018[52] = |(datain[103:100] ^ 1);
  assign w1018[53] = |(datain[99:96] ^ 7);
  assign w1018[54] = |(datain[95:92] ^ 11);
  assign w1018[55] = |(datain[91:88] ^ 4);
  assign w1018[56] = |(datain[87:84] ^ 4);
  assign w1018[57] = |(datain[83:80] ^ 0);
  assign w1018[58] = |(datain[79:76] ^ 11);
  assign w1018[59] = |(datain[75:72] ^ 9);
  assign w1018[60] = |(datain[71:68] ^ 0);
  assign w1018[61] = |(datain[67:64] ^ 3);
  assign w1018[62] = |(datain[63:60] ^ 0);
  assign w1018[63] = |(datain[59:56] ^ 0);
  assign w1018[64] = |(datain[55:52] ^ 11);
  assign w1018[65] = |(datain[51:48] ^ 10);
  assign w1018[66] = |(datain[47:44] ^ 11);
  assign w1018[67] = |(datain[43:40] ^ 3);
  assign w1018[68] = |(datain[39:36] ^ 0);
  assign w1018[69] = |(datain[35:32] ^ 3);
  assign w1018[70] = |(datain[31:28] ^ 12);
  assign w1018[71] = |(datain[27:24] ^ 13);
  assign w1018[72] = |(datain[23:20] ^ 2);
  assign w1018[73] = |(datain[19:16] ^ 1);
  assign comp[1018] = ~(|w1018);
  wire [42-1:0] w1019;
  assign w1019[0] = |(datain[311:308] ^ 11);
  assign w1019[1] = |(datain[307:304] ^ 9);
  assign w1019[2] = |(datain[303:300] ^ 7);
  assign w1019[3] = |(datain[299:296] ^ 10);
  assign w1019[4] = |(datain[295:292] ^ 0);
  assign w1019[5] = |(datain[291:288] ^ 3);
  assign w1019[6] = |(datain[287:284] ^ 11);
  assign w1019[7] = |(datain[283:280] ^ 15);
  assign w1019[8] = |(datain[279:276] ^ 6);
  assign w1019[9] = |(datain[275:272] ^ 3);
  assign w1019[10] = |(datain[271:268] ^ 0);
  assign w1019[11] = |(datain[267:264] ^ 4);
  assign w1019[12] = |(datain[263:260] ^ 8);
  assign w1019[13] = |(datain[259:256] ^ 10);
  assign w1019[14] = |(datain[255:252] ^ 0);
  assign w1019[15] = |(datain[251:248] ^ 4);
  assign w1019[16] = |(datain[247:244] ^ 8);
  assign w1019[17] = |(datain[243:240] ^ 8);
  assign w1019[18] = |(datain[239:236] ^ 0);
  assign w1019[19] = |(datain[235:232] ^ 5);
  assign w1019[20] = |(datain[231:228] ^ 4);
  assign w1019[21] = |(datain[227:224] ^ 7);
  assign w1019[22] = |(datain[223:220] ^ 4);
  assign w1019[23] = |(datain[219:216] ^ 6);
  assign w1019[24] = |(datain[215:212] ^ 14);
  assign w1019[25] = |(datain[211:208] ^ 2);
  assign w1019[26] = |(datain[207:204] ^ 15);
  assign w1019[27] = |(datain[203:200] ^ 8);
  assign w1019[28] = |(datain[199:196] ^ 5);
  assign w1019[29] = |(datain[195:192] ^ 2);
  assign w1019[30] = |(datain[191:188] ^ 11);
  assign w1019[31] = |(datain[187:184] ^ 4);
  assign w1019[32] = |(datain[183:180] ^ 4);
  assign w1019[33] = |(datain[179:176] ^ 0);
  assign w1019[34] = |(datain[175:172] ^ 8);
  assign w1019[35] = |(datain[171:168] ^ 11);
  assign w1019[36] = |(datain[167:164] ^ 1);
  assign w1019[37] = |(datain[163:160] ^ 14);
  assign w1019[38] = |(datain[159:156] ^ 0);
  assign w1019[39] = |(datain[155:152] ^ 15);
  assign w1019[40] = |(datain[151:148] ^ 0);
  assign w1019[41] = |(datain[147:144] ^ 1);
  assign comp[1019] = ~(|w1019);
  wire [74-1:0] w1020;
  assign w1020[0] = |(datain[311:308] ^ 0);
  assign w1020[1] = |(datain[307:304] ^ 2);
  assign w1020[2] = |(datain[303:300] ^ 0);
  assign w1020[3] = |(datain[299:296] ^ 0);
  assign w1020[4] = |(datain[295:292] ^ 8);
  assign w1020[5] = |(datain[291:288] ^ 11);
  assign w1020[6] = |(datain[287:284] ^ 15);
  assign w1020[7] = |(datain[283:280] ^ 0);
  assign w1020[8] = |(datain[279:276] ^ 11);
  assign w1020[9] = |(datain[275:272] ^ 15);
  assign w1020[10] = |(datain[271:268] ^ 3);
  assign w1020[11] = |(datain[267:264] ^ 0);
  assign w1020[12] = |(datain[263:260] ^ 0);
  assign w1020[13] = |(datain[259:256] ^ 1);
  assign w1020[14] = |(datain[255:252] ^ 0);
  assign w1020[15] = |(datain[251:248] ^ 3);
  assign w1020[16] = |(datain[247:244] ^ 15);
  assign w1020[17] = |(datain[243:240] ^ 14);
  assign w1020[18] = |(datain[239:236] ^ 8);
  assign w1020[19] = |(datain[235:232] ^ 10);
  assign w1020[20] = |(datain[231:228] ^ 8);
  assign w1020[21] = |(datain[227:224] ^ 4);
  assign w1020[22] = |(datain[223:220] ^ 13);
  assign w1020[23] = |(datain[219:216] ^ 13);
  assign w1020[24] = |(datain[215:212] ^ 0);
  assign w1020[25] = |(datain[211:208] ^ 6);
  assign w1020[26] = |(datain[207:204] ^ 11);
  assign w1020[27] = |(datain[203:200] ^ 9);
  assign w1020[28] = |(datain[199:196] ^ 10);
  assign w1020[29] = |(datain[195:192] ^ 13);
  assign w1020[30] = |(datain[191:188] ^ 0);
  assign w1020[31] = |(datain[187:184] ^ 5);
  assign w1020[32] = |(datain[183:180] ^ 3);
  assign w1020[33] = |(datain[179:176] ^ 0);
  assign w1020[34] = |(datain[175:172] ^ 0);
  assign w1020[35] = |(datain[171:168] ^ 5);
  assign w1020[36] = |(datain[167:164] ^ 3);
  assign w1020[37] = |(datain[163:160] ^ 12);
  assign w1020[38] = |(datain[159:156] ^ 15);
  assign w1020[39] = |(datain[155:152] ^ 15);
  assign w1020[40] = |(datain[151:148] ^ 7);
  assign w1020[41] = |(datain[147:144] ^ 5);
  assign w1020[42] = |(datain[143:140] ^ 0);
  assign w1020[43] = |(datain[139:136] ^ 2);
  assign w1020[44] = |(datain[135:132] ^ 11);
  assign w1020[45] = |(datain[131:128] ^ 0);
  assign w1020[46] = |(datain[127:124] ^ 0);
  assign w1020[47] = |(datain[123:120] ^ 1);
  assign w1020[48] = |(datain[119:116] ^ 3);
  assign w1020[49] = |(datain[115:112] ^ 12);
  assign w1020[50] = |(datain[111:108] ^ 0);
  assign w1020[51] = |(datain[107:104] ^ 0);
  assign w1020[52] = |(datain[103:100] ^ 7);
  assign w1020[53] = |(datain[99:96] ^ 4);
  assign w1020[54] = |(datain[95:92] ^ 0);
  assign w1020[55] = |(datain[91:88] ^ 2);
  assign w1020[56] = |(datain[87:84] ^ 15);
  assign w1020[57] = |(datain[83:80] ^ 14);
  assign w1020[58] = |(datain[79:76] ^ 12);
  assign w1020[59] = |(datain[75:72] ^ 0);
  assign w1020[60] = |(datain[71:68] ^ 4);
  assign w1020[61] = |(datain[67:64] ^ 7);
  assign w1020[62] = |(datain[63:60] ^ 4);
  assign w1020[63] = |(datain[59:56] ^ 9);
  assign w1020[64] = |(datain[55:52] ^ 8);
  assign w1020[65] = |(datain[51:48] ^ 3);
  assign w1020[66] = |(datain[47:44] ^ 15);
  assign w1020[67] = |(datain[43:40] ^ 9);
  assign w1020[68] = |(datain[39:36] ^ 0);
  assign w1020[69] = |(datain[35:32] ^ 0);
  assign w1020[70] = |(datain[31:28] ^ 7);
  assign w1020[71] = |(datain[27:24] ^ 5);
  assign w1020[72] = |(datain[23:20] ^ 14);
  assign w1020[73] = |(datain[19:16] ^ 11);
  assign comp[1020] = ~(|w1020);
  wire [74-1:0] w1021;
  assign w1021[0] = |(datain[311:308] ^ 12);
  assign w1021[1] = |(datain[307:304] ^ 13);
  assign w1021[2] = |(datain[303:300] ^ 1);
  assign w1021[3] = |(datain[299:296] ^ 3);
  assign w1021[4] = |(datain[295:292] ^ 7);
  assign w1021[5] = |(datain[291:288] ^ 3);
  assign w1021[6] = |(datain[287:284] ^ 0);
  assign w1021[7] = |(datain[283:280] ^ 14);
  assign w1021[8] = |(datain[279:276] ^ 2);
  assign w1021[9] = |(datain[275:272] ^ 14);
  assign w1021[10] = |(datain[271:268] ^ 15);
  assign w1021[11] = |(datain[267:264] ^ 14);
  assign w1021[12] = |(datain[263:260] ^ 0);
  assign w1021[13] = |(datain[259:256] ^ 6);
  assign w1021[14] = |(datain[255:252] ^ 2);
  assign w1021[15] = |(datain[251:248] ^ 0);
  assign w1021[16] = |(datain[247:244] ^ 0);
  assign w1021[17] = |(datain[243:240] ^ 2);
  assign w1021[18] = |(datain[239:236] ^ 2);
  assign w1021[19] = |(datain[235:232] ^ 14);
  assign w1021[20] = |(datain[231:228] ^ 8);
  assign w1021[21] = |(datain[227:224] ^ 0);
  assign w1021[22] = |(datain[223:220] ^ 3);
  assign w1021[23] = |(datain[219:216] ^ 14);
  assign w1021[24] = |(datain[215:212] ^ 2);
  assign w1021[25] = |(datain[211:208] ^ 0);
  assign w1021[26] = |(datain[207:204] ^ 0);
  assign w1021[27] = |(datain[203:200] ^ 2);
  assign w1021[28] = |(datain[199:196] ^ 0);
  assign w1021[29] = |(datain[195:192] ^ 5);
  assign w1021[30] = |(datain[191:188] ^ 7);
  assign w1021[31] = |(datain[187:184] ^ 5);
  assign w1021[32] = |(datain[183:180] ^ 14);
  assign w1021[33] = |(datain[179:176] ^ 6);
  assign w1021[34] = |(datain[175:172] ^ 15);
  assign w1021[35] = |(datain[171:168] ^ 9);
  assign w1021[36] = |(datain[167:164] ^ 12);
  assign w1021[37] = |(datain[163:160] ^ 3);
  assign w1021[38] = |(datain[159:156] ^ 2);
  assign w1021[39] = |(datain[155:152] ^ 14);
  assign w1021[40] = |(datain[151:148] ^ 12);
  assign w1021[41] = |(datain[147:144] ^ 6);
  assign w1021[42] = |(datain[143:140] ^ 0);
  assign w1021[43] = |(datain[139:136] ^ 6);
  assign w1021[44] = |(datain[135:132] ^ 2);
  assign w1021[45] = |(datain[131:128] ^ 0);
  assign w1021[46] = |(datain[127:124] ^ 0);
  assign w1021[47] = |(datain[123:120] ^ 2);
  assign w1021[48] = |(datain[119:116] ^ 0);
  assign w1021[49] = |(datain[115:112] ^ 0);
  assign w1021[50] = |(datain[111:108] ^ 11);
  assign w1021[51] = |(datain[107:104] ^ 8);
  assign w1021[52] = |(datain[103:100] ^ 0);
  assign w1021[53] = |(datain[99:96] ^ 1);
  assign w1021[54] = |(datain[95:92] ^ 0);
  assign w1021[55] = |(datain[91:88] ^ 3);
  assign w1021[56] = |(datain[87:84] ^ 11);
  assign w1021[57] = |(datain[83:80] ^ 11);
  assign w1021[58] = |(datain[79:76] ^ 0);
  assign w1021[59] = |(datain[75:72] ^ 0);
  assign w1021[60] = |(datain[71:68] ^ 7);
  assign w1021[61] = |(datain[67:64] ^ 12);
  assign w1021[62] = |(datain[63:60] ^ 11);
  assign w1021[63] = |(datain[59:56] ^ 14);
  assign w1021[64] = |(datain[55:52] ^ 0);
  assign w1021[65] = |(datain[51:48] ^ 10);
  assign w1021[66] = |(datain[47:44] ^ 0);
  assign w1021[67] = |(datain[43:40] ^ 7);
  assign w1021[68] = |(datain[39:36] ^ 12);
  assign w1021[69] = |(datain[35:32] ^ 13);
  assign w1021[70] = |(datain[31:28] ^ 1);
  assign w1021[71] = |(datain[27:24] ^ 3);
  assign w1021[72] = |(datain[23:20] ^ 7);
  assign w1021[73] = |(datain[19:16] ^ 3);
  assign comp[1021] = ~(|w1021);
  wire [66-1:0] w1022;
  assign w1022[0] = |(datain[311:308] ^ 0);
  assign w1022[1] = |(datain[307:304] ^ 1);
  assign w1022[2] = |(datain[303:300] ^ 8);
  assign w1022[3] = |(datain[299:296] ^ 11);
  assign w1022[4] = |(datain[295:292] ^ 0);
  assign w1022[5] = |(datain[291:288] ^ 5);
  assign w1022[6] = |(datain[287:284] ^ 2);
  assign w1022[7] = |(datain[283:280] ^ 13);
  assign w1022[8] = |(datain[279:276] ^ 0);
  assign w1022[9] = |(datain[275:272] ^ 2);
  assign w1022[10] = |(datain[271:268] ^ 0);
  assign w1022[11] = |(datain[267:264] ^ 0);
  assign w1022[12] = |(datain[263:260] ^ 8);
  assign w1022[13] = |(datain[259:256] ^ 11);
  assign w1022[14] = |(datain[255:252] ^ 15);
  assign w1022[15] = |(datain[251:248] ^ 0);
  assign w1022[16] = |(datain[247:244] ^ 8);
  assign w1022[17] = |(datain[243:240] ^ 10);
  assign w1022[18] = |(datain[239:236] ^ 8);
  assign w1022[19] = |(datain[235:232] ^ 4);
  assign w1022[20] = |(datain[231:228] ^ 9);
  assign w1022[21] = |(datain[227:224] ^ 9);
  assign w1022[22] = |(datain[223:220] ^ 0);
  assign w1022[23] = |(datain[219:216] ^ 4);
  assign w1022[24] = |(datain[215:212] ^ 11);
  assign w1022[25] = |(datain[211:208] ^ 11);
  assign w1022[26] = |(datain[207:204] ^ 2);
  assign w1022[27] = |(datain[203:200] ^ 8);
  assign w1022[28] = |(datain[199:196] ^ 0);
  assign w1022[29] = |(datain[195:192] ^ 1);
  assign w1022[30] = |(datain[191:188] ^ 0);
  assign w1022[31] = |(datain[187:184] ^ 3);
  assign w1022[32] = |(datain[183:180] ^ 13);
  assign w1022[33] = |(datain[179:176] ^ 14);
  assign w1022[34] = |(datain[175:172] ^ 11);
  assign w1022[35] = |(datain[171:168] ^ 9);
  assign w1022[36] = |(datain[167:164] ^ 7);
  assign w1022[37] = |(datain[163:160] ^ 1);
  assign w1022[38] = |(datain[159:156] ^ 0);
  assign w1022[39] = |(datain[155:152] ^ 3);
  assign w1022[40] = |(datain[151:148] ^ 8);
  assign w1022[41] = |(datain[147:144] ^ 10);
  assign w1022[42] = |(datain[143:140] ^ 2);
  assign w1022[43] = |(datain[139:136] ^ 7);
  assign w1022[44] = |(datain[135:132] ^ 3);
  assign w1022[45] = |(datain[131:128] ^ 2);
  assign w1022[46] = |(datain[127:124] ^ 14);
  assign w1022[47] = |(datain[123:120] ^ 0);
  assign w1022[48] = |(datain[119:116] ^ 8);
  assign w1022[49] = |(datain[115:112] ^ 8);
  assign w1022[50] = |(datain[111:108] ^ 2);
  assign w1022[51] = |(datain[107:104] ^ 7);
  assign w1022[52] = |(datain[103:100] ^ 4);
  assign w1022[53] = |(datain[99:96] ^ 3);
  assign w1022[54] = |(datain[95:92] ^ 4);
  assign w1022[55] = |(datain[91:88] ^ 9);
  assign w1022[56] = |(datain[87:84] ^ 8);
  assign w1022[57] = |(datain[83:80] ^ 3);
  assign w1022[58] = |(datain[79:76] ^ 15);
  assign w1022[59] = |(datain[75:72] ^ 9);
  assign w1022[60] = |(datain[71:68] ^ 0);
  assign w1022[61] = |(datain[67:64] ^ 0);
  assign w1022[62] = |(datain[63:60] ^ 7);
  assign w1022[63] = |(datain[59:56] ^ 5);
  assign w1022[64] = |(datain[55:52] ^ 15);
  assign w1022[65] = |(datain[51:48] ^ 3);
  assign comp[1022] = ~(|w1022);
  wire [73-1:0] w1023;
  assign w1023[0] = |(datain[311:308] ^ 11);
  assign w1023[1] = |(datain[307:304] ^ 9);
  assign w1023[2] = |(datain[303:300] ^ 6);
  assign w1023[3] = |(datain[299:296] ^ 8);
  assign w1023[4] = |(datain[295:292] ^ 0);
  assign w1023[5] = |(datain[291:288] ^ 3);
  assign w1023[6] = |(datain[287:284] ^ 11);
  assign w1023[7] = |(datain[283:280] ^ 4);
  assign w1023[8] = |(datain[279:276] ^ 4);
  assign w1023[9] = |(datain[275:272] ^ 0);
  assign w1023[10] = |(datain[271:268] ^ 12);
  assign w1023[11] = |(datain[267:264] ^ 12);
  assign w1023[12] = |(datain[263:260] ^ 3);
  assign w1023[13] = |(datain[259:256] ^ 3);
  assign w1023[14] = |(datain[255:252] ^ 12);
  assign w1023[15] = |(datain[251:248] ^ 9);
  assign w1023[16] = |(datain[247:244] ^ 8);
  assign w1023[17] = |(datain[243:240] ^ 1);
  assign w1023[18] = |(datain[239:236] ^ 14);
  assign w1023[19] = |(datain[235:232] ^ 15);
  assign w1023[20] = |(datain[231:228] ^ 15);
  assign w1023[21] = |(datain[227:224] ^ 15);
  assign w1023[22] = |(datain[223:220] ^ 0);
  assign w1023[23] = |(datain[219:216] ^ 0);
  assign w1023[24] = |(datain[215:212] ^ 8);
  assign w1023[25] = |(datain[211:208] ^ 11);
  assign w1023[26] = |(datain[207:204] ^ 13);
  assign w1023[27] = |(datain[203:200] ^ 7);
  assign w1023[28] = |(datain[199:196] ^ 11);
  assign w1023[29] = |(datain[195:192] ^ 8);
  assign w1023[30] = |(datain[191:188] ^ 0);
  assign w1023[31] = |(datain[187:184] ^ 0);
  assign w1023[32] = |(datain[183:180] ^ 4);
  assign w1023[33] = |(datain[179:176] ^ 2);
  assign w1023[34] = |(datain[175:172] ^ 12);
  assign w1023[35] = |(datain[171:168] ^ 12);
  assign w1023[36] = |(datain[167:164] ^ 11);
  assign w1023[37] = |(datain[163:160] ^ 10);
  assign w1023[38] = |(datain[159:156] ^ 7);
  assign w1023[39] = |(datain[155:152] ^ 2);
  assign w1023[40] = |(datain[151:148] ^ 0);
  assign w1023[41] = |(datain[147:144] ^ 3);
  assign w1023[42] = |(datain[143:140] ^ 11);
  assign w1023[43] = |(datain[139:136] ^ 9);
  assign w1023[44] = |(datain[135:132] ^ 0);
  assign w1023[45] = |(datain[131:128] ^ 2);
  assign w1023[46] = |(datain[127:124] ^ 0);
  assign w1023[47] = |(datain[123:120] ^ 0);
  assign w1023[48] = |(datain[119:116] ^ 11);
  assign w1023[49] = |(datain[115:112] ^ 4);
  assign w1023[50] = |(datain[111:108] ^ 4);
  assign w1023[51] = |(datain[107:104] ^ 0);
  assign w1023[52] = |(datain[103:100] ^ 12);
  assign w1023[53] = |(datain[99:96] ^ 12);
  assign w1023[54] = |(datain[95:92] ^ 14);
  assign w1023[55] = |(datain[91:88] ^ 8);
  assign w1023[56] = |(datain[87:84] ^ 5);
  assign w1023[57] = |(datain[83:80] ^ 1);
  assign w1023[58] = |(datain[79:76] ^ 0);
  assign w1023[59] = |(datain[75:72] ^ 0);
  assign w1023[60] = |(datain[71:68] ^ 11);
  assign w1023[61] = |(datain[67:64] ^ 4);
  assign w1023[62] = |(datain[63:60] ^ 3);
  assign w1023[63] = |(datain[59:56] ^ 14);
  assign w1023[64] = |(datain[55:52] ^ 12);
  assign w1023[65] = |(datain[51:48] ^ 12);
  assign w1023[66] = |(datain[47:44] ^ 11);
  assign w1023[67] = |(datain[43:40] ^ 10);
  assign w1023[68] = |(datain[39:36] ^ 7);
  assign w1023[69] = |(datain[35:32] ^ 11);
  assign w1023[70] = |(datain[31:28] ^ 0);
  assign w1023[71] = |(datain[27:24] ^ 3);
  assign w1023[72] = |(datain[23:20] ^ 14);
  assign w1023[73] = |(datain[19:16] ^ 8);
  assign comp[1023] = ~(|w1023);
  wire [11-1:0] dout_wr;

  always @(posedge clk) begin
    if(rst) begin
      dout <= 0;
    end else begin
      dout <= dout_wr;
    end
  end

generate
  genvar n;
  for(n=0;n<1024;n=n+1)
  begin: shifters
    assign dout_wr = comp[n] ? n: {11{1'bz}};
  end
endgenerate

endmodule

